magic
tech sky130A
magscale 1 2
timestamp 1639277212
<< checkpaint >>
rect -12658 -11586 596582 715522
<< locali >>
rect 252569 486659 252603 486965
rect 253857 486251 253891 486965
rect 257905 486319 257939 487033
rect 261861 486387 261895 486965
rect 264437 486455 264471 486965
rect 265725 486523 265759 486965
rect 345305 486115 345339 487577
rect 355609 486047 355643 487509
rect 359473 485979 359507 487509
rect 363429 485911 363463 487509
rect 367293 485843 367327 487509
rect 265449 335971 265483 336481
rect 351929 336311 351963 336549
rect 364165 336549 364257 336583
rect 352021 336175 352055 336345
rect 351871 336141 352055 336175
rect 353309 336107 353343 336277
rect 362693 335631 362727 336005
rect 364165 335767 364199 336549
rect 382197 335903 382231 336753
rect 380725 335835 380759 335869
rect 380633 335801 380759 335835
rect 380633 335767 380667 335801
rect 370881 335495 370915 335597
rect 377505 335563 377539 335733
rect 379379 335665 379471 335699
rect 371893 335427 371927 335529
rect 379437 335427 379471 335665
rect 380725 335359 380759 335733
rect 295533 323595 295567 326485
rect 249717 6919 249751 7769
rect 249935 7633 250085 7667
rect 234537 4879 234571 4913
rect 234537 4845 234813 4879
rect 243461 4845 243679 4879
rect 231961 4267 231995 4777
rect 243461 4267 243495 4845
rect 243645 4811 243679 4845
rect 244841 4811 244875 4913
rect 244841 4777 245025 4811
rect 243553 4267 243587 4777
rect 240149 4199 240183 4233
rect 240149 4165 240333 4199
rect 241529 3587 241563 4097
rect 256709 3383 256743 3553
rect 290657 3111 290691 3349
rect 299581 3179 299615 3349
rect 301053 3247 301087 3689
rect 305377 3315 305411 4097
rect 330585 3723 330619 3893
rect 306481 3587 306515 3689
rect 331689 3587 331723 4097
rect 333713 4097 334081 4131
rect 333713 3859 333747 4097
rect 333989 3995 334023 4029
rect 333989 3961 334265 3995
rect 336749 3961 336933 3995
rect 336749 3927 336783 3961
rect 324513 3315 324547 3417
rect 298017 2839 298051 3077
rect 301605 2771 301639 3281
rect 333621 2771 333655 3689
rect 334173 3519 334207 3893
rect 334265 3315 334299 3485
rect 334357 2907 334391 3281
rect 427093 2907 427127 3689
rect 429761 2975 429795 3757
rect 440433 3043 440467 3757
rect 446321 3077 446505 3111
rect 446321 3043 446355 3077
rect 436845 2907 436879 3009
rect 436695 2873 436879 2907
rect 334299 2805 334541 2839
rect 427035 2805 427277 2839
<< viali >>
rect 345305 487577 345339 487611
rect 257905 487033 257939 487067
rect 252569 486965 252603 486999
rect 252569 486625 252603 486659
rect 253857 486965 253891 486999
rect 261861 486965 261895 486999
rect 264437 486965 264471 486999
rect 265725 486965 265759 486999
rect 265725 486489 265759 486523
rect 264437 486421 264471 486455
rect 261861 486353 261895 486387
rect 257905 486285 257939 486319
rect 253857 486217 253891 486251
rect 345305 486081 345339 486115
rect 355609 487509 355643 487543
rect 355609 486013 355643 486047
rect 359473 487509 359507 487543
rect 359473 485945 359507 485979
rect 363429 487509 363463 487543
rect 363429 485877 363463 485911
rect 367293 487509 367327 487543
rect 367293 485809 367327 485843
rect 382197 336753 382231 336787
rect 351929 336549 351963 336583
rect 265449 336481 265483 336515
rect 364257 336549 364291 336583
rect 351929 336277 351963 336311
rect 352021 336345 352055 336379
rect 351837 336141 351871 336175
rect 353309 336277 353343 336311
rect 353309 336073 353343 336107
rect 265449 335937 265483 335971
rect 362693 336005 362727 336039
rect 380725 335869 380759 335903
rect 382197 335869 382231 335903
rect 364165 335733 364199 335767
rect 377505 335733 377539 335767
rect 380633 335733 380667 335767
rect 380725 335733 380759 335767
rect 362693 335597 362727 335631
rect 370881 335597 370915 335631
rect 379345 335665 379379 335699
rect 370881 335461 370915 335495
rect 371893 335529 371927 335563
rect 377505 335529 377539 335563
rect 371893 335393 371927 335427
rect 379437 335393 379471 335427
rect 380725 335325 380759 335359
rect 295533 326485 295567 326519
rect 295533 323561 295567 323595
rect 249717 7769 249751 7803
rect 249901 7633 249935 7667
rect 250085 7633 250119 7667
rect 249717 6885 249751 6919
rect 234537 4913 234571 4947
rect 244841 4913 244875 4947
rect 234813 4845 234847 4879
rect 231961 4777 231995 4811
rect 231961 4233 231995 4267
rect 240149 4233 240183 4267
rect 243461 4233 243495 4267
rect 243553 4777 243587 4811
rect 243645 4777 243679 4811
rect 245025 4777 245059 4811
rect 243553 4233 243587 4267
rect 240333 4165 240367 4199
rect 241529 4097 241563 4131
rect 305377 4097 305411 4131
rect 301053 3689 301087 3723
rect 241529 3553 241563 3587
rect 256709 3553 256743 3587
rect 256709 3349 256743 3383
rect 290657 3349 290691 3383
rect 299581 3349 299615 3383
rect 331689 4097 331723 4131
rect 330585 3893 330619 3927
rect 306481 3689 306515 3723
rect 330585 3689 330619 3723
rect 306481 3553 306515 3587
rect 334081 4097 334115 4131
rect 333989 4029 334023 4063
rect 334265 3961 334299 3995
rect 336933 3961 336967 3995
rect 333713 3825 333747 3859
rect 334173 3893 334207 3927
rect 336749 3893 336783 3927
rect 331689 3553 331723 3587
rect 333621 3689 333655 3723
rect 301053 3213 301087 3247
rect 301605 3281 301639 3315
rect 305377 3281 305411 3315
rect 324513 3417 324547 3451
rect 324513 3281 324547 3315
rect 299581 3145 299615 3179
rect 290657 3077 290691 3111
rect 298017 3077 298051 3111
rect 298017 2805 298051 2839
rect 301605 2737 301639 2771
rect 429761 3757 429795 3791
rect 427093 3689 427127 3723
rect 334173 3485 334207 3519
rect 334265 3485 334299 3519
rect 334265 3281 334299 3315
rect 334357 3281 334391 3315
rect 334357 2873 334391 2907
rect 440433 3757 440467 3791
rect 429761 2941 429795 2975
rect 436845 3009 436879 3043
rect 440433 3009 440467 3043
rect 446505 3077 446539 3111
rect 446321 3009 446355 3043
rect 427093 2873 427127 2907
rect 436661 2873 436695 2907
rect 334265 2805 334299 2839
rect 334541 2805 334575 2839
rect 427001 2805 427035 2839
rect 427277 2805 427311 2839
rect 333621 2737 333655 2771
<< metal1 >>
rect 170306 700952 170312 701004
rect 170364 700992 170370 701004
rect 316034 700992 316040 701004
rect 170364 700964 316040 700992
rect 170364 700952 170370 700964
rect 316034 700952 316040 700964
rect 316092 700952 316098 701004
rect 154114 700884 154120 700936
rect 154172 700924 154178 700936
rect 312538 700924 312544 700936
rect 154172 700896 312544 700924
rect 154172 700884 154178 700896
rect 312538 700884 312544 700896
rect 312596 700884 312602 700936
rect 299382 700816 299388 700868
rect 299440 700856 299446 700868
rect 462314 700856 462320 700868
rect 299440 700828 462320 700856
rect 299440 700816 299446 700828
rect 462314 700816 462320 700828
rect 462372 700816 462378 700868
rect 300762 700748 300768 700800
rect 300820 700788 300826 700800
rect 478506 700788 478512 700800
rect 300820 700760 478512 700788
rect 300820 700748 300826 700760
rect 478506 700748 478512 700760
rect 478564 700748 478570 700800
rect 137830 700680 137836 700732
rect 137888 700720 137894 700732
rect 317414 700720 317420 700732
rect 137888 700692 317420 700720
rect 137888 700680 137894 700692
rect 317414 700680 317420 700692
rect 317472 700680 317478 700732
rect 298002 700612 298008 700664
rect 298060 700652 298066 700664
rect 494790 700652 494796 700664
rect 298060 700624 494796 700652
rect 298060 700612 298066 700624
rect 494790 700612 494796 700624
rect 494848 700612 494854 700664
rect 105446 700544 105452 700596
rect 105504 700584 105510 700596
rect 320174 700584 320180 700596
rect 105504 700556 320180 700584
rect 105504 700544 105510 700556
rect 320174 700544 320180 700556
rect 320232 700544 320238 700596
rect 89162 700476 89168 700528
rect 89220 700516 89226 700528
rect 315298 700516 315304 700528
rect 89220 700488 315304 700516
rect 89220 700476 89226 700488
rect 315298 700476 315304 700488
rect 315356 700476 315362 700528
rect 295242 700408 295248 700460
rect 295300 700448 295306 700460
rect 527174 700448 527180 700460
rect 295300 700420 527180 700448
rect 295300 700408 295306 700420
rect 527174 700408 527180 700420
rect 527232 700408 527238 700460
rect 296622 700340 296628 700392
rect 296680 700380 296686 700392
rect 543458 700380 543464 700392
rect 296680 700352 543464 700380
rect 296680 700340 296686 700352
rect 543458 700340 543464 700352
rect 543516 700340 543522 700392
rect 72970 700272 72976 700324
rect 73028 700312 73034 700324
rect 321554 700312 321560 700324
rect 73028 700284 321560 700312
rect 73028 700272 73034 700284
rect 321554 700272 321560 700284
rect 321612 700272 321618 700324
rect 302142 700204 302148 700256
rect 302200 700244 302206 700256
rect 429838 700244 429844 700256
rect 302200 700216 429844 700244
rect 302200 700204 302206 700216
rect 429838 700204 429844 700216
rect 429896 700204 429902 700256
rect 202782 700136 202788 700188
rect 202840 700176 202846 700188
rect 313274 700176 313280 700188
rect 202840 700148 313280 700176
rect 202840 700136 202846 700148
rect 313274 700136 313280 700148
rect 313332 700136 313338 700188
rect 304902 700068 304908 700120
rect 304960 700108 304966 700120
rect 413646 700108 413652 700120
rect 304960 700080 413652 700108
rect 304960 700068 304966 700080
rect 413646 700068 413652 700080
rect 413704 700068 413710 700120
rect 303522 700000 303528 700052
rect 303580 700040 303586 700052
rect 397454 700040 397460 700052
rect 303580 700012 397460 700040
rect 303580 700000 303586 700012
rect 397454 700000 397460 700012
rect 397512 700000 397518 700052
rect 235166 699932 235172 699984
rect 235224 699972 235230 699984
rect 311986 699972 311992 699984
rect 235224 699944 311992 699972
rect 235224 699932 235230 699944
rect 311986 699932 311992 699944
rect 312044 699932 312050 699984
rect 306282 699864 306288 699916
rect 306340 699904 306346 699916
rect 364978 699904 364984 699916
rect 306340 699876 364984 699904
rect 306340 699864 306346 699876
rect 364978 699864 364984 699876
rect 365036 699864 365042 699916
rect 267642 699796 267648 699848
rect 267700 699836 267706 699848
rect 310514 699836 310520 699848
rect 267700 699808 310520 699836
rect 267700 699796 267706 699808
rect 310514 699796 310520 699808
rect 310572 699796 310578 699848
rect 307662 699728 307668 699780
rect 307720 699768 307726 699780
rect 332502 699768 332508 699780
rect 307720 699740 332508 699768
rect 307720 699728 307726 699740
rect 332502 699728 332508 699740
rect 332560 699728 332566 699780
rect 300118 699660 300124 699712
rect 300176 699700 300182 699712
rect 309134 699700 309140 699712
rect 300176 699672 309140 699700
rect 300176 699660 300182 699672
rect 309134 699660 309140 699672
rect 309192 699660 309198 699712
rect 292482 696940 292488 696992
rect 292540 696980 292546 696992
rect 580166 696980 580172 696992
rect 292540 696952 580172 696980
rect 292540 696940 292546 696952
rect 580166 696940 580172 696952
rect 580224 696940 580230 696992
rect 292390 683204 292396 683256
rect 292448 683244 292454 683256
rect 580166 683244 580172 683256
rect 292448 683216 580172 683244
rect 292448 683204 292454 683216
rect 580166 683204 580172 683216
rect 580224 683204 580230 683256
rect 3418 683136 3424 683188
rect 3476 683176 3482 683188
rect 328454 683176 328460 683188
rect 3476 683148 328460 683176
rect 3476 683136 3482 683148
rect 328454 683136 328460 683148
rect 328512 683136 328518 683188
rect 291102 670760 291108 670812
rect 291160 670800 291166 670812
rect 580166 670800 580172 670812
rect 291160 670772 580172 670800
rect 291160 670760 291166 670772
rect 580166 670760 580172 670772
rect 580224 670760 580230 670812
rect 3510 670692 3516 670744
rect 3568 670732 3574 670744
rect 323578 670732 323584 670744
rect 3568 670704 323584 670732
rect 3568 670692 3574 670704
rect 323578 670692 323584 670704
rect 323636 670692 323642 670744
rect 3418 656888 3424 656940
rect 3476 656928 3482 656940
rect 329834 656928 329840 656940
rect 3476 656900 329840 656928
rect 3476 656888 3482 656900
rect 329834 656888 329840 656900
rect 329892 656888 329898 656940
rect 288342 643084 288348 643136
rect 288400 643124 288406 643136
rect 580166 643124 580172 643136
rect 288400 643096 580172 643124
rect 288400 643084 288406 643096
rect 580166 643084 580172 643096
rect 580224 643084 580230 643136
rect 3418 632068 3424 632120
rect 3476 632108 3482 632120
rect 332594 632108 332600 632120
rect 3476 632080 332600 632108
rect 3476 632068 3482 632080
rect 332594 632068 332600 632080
rect 332652 632068 332658 632120
rect 289722 630640 289728 630692
rect 289780 630680 289786 630692
rect 580166 630680 580172 630692
rect 289780 630652 580172 630680
rect 289780 630640 289786 630652
rect 580166 630640 580172 630652
rect 580224 630640 580230 630692
rect 3142 618264 3148 618316
rect 3200 618304 3206 618316
rect 327718 618304 327724 618316
rect 3200 618276 327724 618304
rect 3200 618264 3206 618276
rect 327718 618264 327724 618276
rect 327776 618264 327782 618316
rect 286962 616836 286968 616888
rect 287020 616876 287026 616888
rect 580166 616876 580172 616888
rect 287020 616848 580172 616876
rect 287020 616836 287026 616848
rect 580166 616836 580172 616848
rect 580224 616836 580230 616888
rect 3234 605820 3240 605872
rect 3292 605860 3298 605872
rect 332686 605860 332692 605872
rect 3292 605832 332692 605860
rect 3292 605820 3298 605832
rect 332686 605820 332692 605832
rect 332744 605820 332750 605872
rect 284110 590656 284116 590708
rect 284168 590696 284174 590708
rect 579798 590696 579804 590708
rect 284168 590668 579804 590696
rect 284168 590656 284174 590668
rect 579798 590656 579804 590668
rect 579856 590656 579862 590708
rect 3326 579640 3332 579692
rect 3384 579680 3390 579692
rect 335354 579680 335360 579692
rect 3384 579652 335360 579680
rect 3384 579640 3390 579652
rect 335354 579640 335360 579652
rect 335412 579640 335418 579692
rect 285582 576852 285588 576904
rect 285640 576892 285646 576904
rect 580166 576892 580172 576904
rect 285640 576864 580172 576892
rect 285640 576852 285646 576864
rect 580166 576852 580172 576864
rect 580224 576852 580230 576904
rect 3418 565836 3424 565888
rect 3476 565876 3482 565888
rect 331858 565876 331864 565888
rect 3476 565848 331864 565876
rect 3476 565836 3482 565848
rect 331858 565836 331864 565848
rect 331916 565836 331922 565888
rect 282822 563048 282828 563100
rect 282880 563088 282886 563100
rect 579798 563088 579804 563100
rect 282880 563060 579804 563088
rect 282880 563048 282886 563060
rect 579798 563048 579804 563060
rect 579856 563048 579862 563100
rect 3418 553392 3424 553444
rect 3476 553432 3482 553444
rect 336734 553432 336740 553444
rect 3476 553404 336740 553432
rect 3476 553392 3482 553404
rect 336734 553392 336740 553404
rect 336792 553392 336798 553444
rect 280062 536800 280068 536852
rect 280120 536840 280126 536852
rect 580166 536840 580172 536852
rect 280120 536812 580172 536840
rect 280120 536800 280126 536812
rect 580166 536800 580172 536812
rect 580224 536800 580230 536852
rect 3418 527144 3424 527196
rect 3476 527184 3482 527196
rect 339494 527184 339500 527196
rect 3476 527156 339500 527184
rect 3476 527144 3482 527156
rect 339494 527144 339500 527156
rect 339552 527144 339558 527196
rect 281442 524424 281448 524476
rect 281500 524464 281506 524476
rect 580166 524464 580172 524476
rect 281500 524436 580172 524464
rect 281500 524424 281506 524436
rect 580166 524424 580172 524436
rect 580224 524424 580230 524476
rect 3418 514768 3424 514820
rect 3476 514808 3482 514820
rect 334618 514808 334624 514820
rect 3476 514780 334624 514808
rect 3476 514768 3482 514780
rect 334618 514768 334624 514780
rect 334676 514768 334682 514820
rect 278682 510620 278688 510672
rect 278740 510660 278746 510672
rect 580166 510660 580172 510672
rect 278740 510632 580172 510660
rect 278740 510620 278746 510632
rect 580166 510620 580172 510632
rect 580224 510620 580230 510672
rect 3050 500964 3056 501016
rect 3108 501004 3114 501016
rect 340874 501004 340880 501016
rect 3108 500976 340880 501004
rect 3108 500964 3114 500976
rect 340874 500964 340880 500976
rect 340932 500964 340938 501016
rect 285122 491240 285128 491292
rect 285180 491280 285186 491292
rect 285582 491280 285588 491292
rect 285180 491252 285588 491280
rect 285180 491240 285186 491252
rect 285582 491240 285588 491252
rect 285640 491240 285646 491292
rect 286410 491240 286416 491292
rect 286468 491280 286474 491292
rect 286962 491280 286968 491292
rect 286468 491252 286968 491280
rect 286468 491240 286474 491252
rect 286962 491240 286968 491252
rect 287020 491240 287026 491292
rect 287698 491240 287704 491292
rect 287756 491280 287762 491292
rect 288342 491280 288348 491292
rect 287756 491252 288348 491280
rect 287756 491240 287762 491252
rect 288342 491240 288348 491252
rect 288400 491240 288406 491292
rect 288986 491240 288992 491292
rect 289044 491280 289050 491292
rect 289722 491280 289728 491292
rect 289044 491252 289728 491280
rect 289044 491240 289050 491252
rect 289722 491240 289728 491252
rect 289780 491240 289786 491292
rect 290274 491240 290280 491292
rect 290332 491280 290338 491292
rect 291102 491280 291108 491292
rect 290332 491252 291108 491280
rect 290332 491240 290338 491252
rect 291102 491240 291108 491252
rect 291160 491240 291166 491292
rect 291562 491240 291568 491292
rect 291620 491280 291626 491292
rect 292482 491280 292488 491292
rect 291620 491252 292488 491280
rect 291620 491240 291626 491252
rect 292482 491240 292488 491252
rect 292540 491240 292546 491292
rect 305822 491240 305828 491292
rect 305880 491280 305886 491292
rect 306282 491280 306288 491292
rect 305880 491252 306288 491280
rect 305880 491240 305886 491252
rect 306282 491240 306288 491252
rect 306340 491240 306346 491292
rect 307110 491240 307116 491292
rect 307168 491280 307174 491292
rect 307662 491280 307668 491292
rect 307168 491252 307668 491280
rect 307168 491240 307174 491252
rect 307662 491240 307668 491252
rect 307720 491240 307726 491292
rect 327718 491240 327724 491292
rect 327776 491280 327782 491292
rect 334894 491280 334900 491292
rect 327776 491252 334900 491280
rect 327776 491240 327782 491252
rect 334894 491240 334900 491252
rect 334952 491240 334958 491292
rect 284202 491172 284208 491224
rect 284260 491212 284266 491224
rect 311894 491212 311900 491224
rect 284260 491184 311900 491212
rect 284260 491172 284266 491184
rect 311894 491172 311900 491184
rect 311952 491172 311958 491224
rect 312538 491172 312544 491224
rect 312596 491212 312602 491224
rect 319346 491212 319352 491224
rect 312596 491184 319352 491212
rect 312596 491172 312602 491184
rect 319346 491172 319352 491184
rect 319404 491172 319410 491224
rect 319438 491172 319444 491224
rect 319496 491212 319502 491224
rect 327166 491212 327172 491224
rect 319496 491184 327172 491212
rect 319496 491172 319502 491184
rect 327166 491172 327172 491184
rect 327224 491172 327230 491224
rect 331858 491172 331864 491224
rect 331916 491212 331922 491224
rect 338758 491212 338764 491224
rect 331916 491184 338764 491212
rect 331916 491172 331922 491184
rect 338758 491172 338764 491184
rect 338816 491172 338822 491224
rect 308398 491104 308404 491156
rect 308456 491144 308462 491156
rect 347774 491144 347780 491156
rect 308456 491116 347780 491144
rect 308456 491104 308462 491116
rect 347774 491104 347780 491116
rect 347832 491104 347838 491156
rect 219342 491036 219348 491088
rect 219400 491076 219406 491088
rect 315206 491076 315212 491088
rect 219400 491048 315212 491076
rect 219400 491036 219406 491048
rect 315206 491036 315212 491048
rect 315264 491036 315270 491088
rect 315298 491036 315304 491088
rect 315356 491076 315362 491088
rect 323302 491076 323308 491088
rect 315356 491048 323308 491076
rect 315356 491036 315362 491048
rect 323302 491036 323308 491048
rect 323360 491036 323366 491088
rect 323578 491036 323584 491088
rect 323636 491076 323642 491088
rect 331214 491076 331220 491088
rect 323636 491048 331220 491076
rect 323636 491036 323642 491048
rect 331214 491036 331220 491048
rect 331272 491036 331278 491088
rect 334618 491036 334624 491088
rect 334676 491076 334682 491088
rect 342714 491076 342720 491088
rect 334676 491048 342720 491076
rect 334676 491036 334682 491048
rect 342714 491036 342720 491048
rect 342772 491036 342778 491088
rect 273162 490968 273168 491020
rect 273220 491008 273226 491020
rect 385954 491008 385960 491020
rect 273220 490980 385960 491008
rect 273220 490968 273226 490980
rect 385954 490968 385960 490980
rect 386012 490968 386018 491020
rect 271782 490900 271788 490952
rect 271840 490940 271846 490952
rect 386046 490940 386052 490952
rect 271840 490912 386052 490940
rect 271840 490900 271846 490912
rect 386046 490900 386052 490912
rect 386104 490900 386110 490952
rect 7926 490832 7932 490884
rect 7984 490872 7990 490884
rect 346578 490872 346584 490884
rect 7984 490844 346584 490872
rect 7984 490832 7990 490844
rect 346578 490832 346584 490844
rect 346636 490832 346642 490884
rect 5442 490764 5448 490816
rect 5500 490804 5506 490816
rect 347958 490804 347964 490816
rect 5500 490776 347964 490804
rect 5500 490764 5506 490776
rect 347958 490764 347964 490776
rect 348016 490764 348022 490816
rect 5350 490696 5356 490748
rect 5408 490736 5414 490748
rect 349154 490736 349160 490748
rect 5408 490708 349160 490736
rect 5408 490696 5414 490708
rect 349154 490696 349160 490708
rect 349212 490696 349218 490748
rect 5258 490628 5264 490680
rect 5316 490668 5322 490680
rect 351914 490668 351920 490680
rect 5316 490640 351920 490668
rect 5316 490628 5322 490640
rect 351914 490628 351920 490640
rect 351972 490628 351978 490680
rect 3326 490560 3332 490612
rect 3384 490600 3390 490612
rect 350534 490600 350540 490612
rect 3384 490572 350540 490600
rect 3384 490560 3390 490572
rect 350534 490560 350540 490572
rect 350592 490560 350598 490612
rect 4062 490492 4068 490544
rect 4120 490532 4126 490544
rect 354306 490532 354312 490544
rect 4120 490504 354312 490532
rect 4120 490492 4126 490504
rect 354306 490492 354312 490504
rect 354364 490492 354370 490544
rect 3970 490424 3976 490476
rect 4028 490464 4034 490476
rect 353294 490464 353300 490476
rect 4028 490436 353300 490464
rect 4028 490424 4034 490436
rect 353294 490424 353300 490436
rect 353352 490424 353358 490476
rect 6546 490356 6552 490408
rect 6604 490396 6610 490408
rect 356882 490396 356888 490408
rect 6604 490368 356888 490396
rect 6604 490356 6610 490368
rect 356882 490356 356888 490368
rect 356940 490356 356946 490408
rect 3878 490288 3884 490340
rect 3936 490328 3942 490340
rect 358170 490328 358176 490340
rect 3936 490300 358176 490328
rect 3936 490288 3942 490300
rect 358170 490288 358176 490300
rect 358228 490288 358234 490340
rect 6454 490220 6460 490272
rect 6512 490260 6518 490272
rect 360746 490260 360752 490272
rect 6512 490232 360752 490260
rect 6512 490220 6518 490232
rect 360746 490220 360752 490232
rect 360804 490220 360810 490272
rect 3786 490152 3792 490204
rect 3844 490192 3850 490204
rect 362126 490192 362132 490204
rect 3844 490164 362132 490192
rect 3844 490152 3850 490164
rect 362126 490152 362132 490164
rect 362184 490152 362190 490204
rect 6362 490084 6368 490136
rect 6420 490124 6426 490136
rect 364702 490124 364708 490136
rect 6420 490096 364708 490124
rect 6420 490084 6426 490096
rect 364702 490084 364708 490096
rect 364760 490084 364766 490136
rect 3602 490016 3608 490068
rect 3660 490056 3666 490068
rect 365990 490056 365996 490068
rect 3660 490028 365996 490056
rect 3660 490016 3666 490028
rect 365990 490016 365996 490028
rect 366048 490016 366054 490068
rect 6270 489948 6276 490000
rect 6328 489988 6334 490000
rect 368566 489988 368572 490000
rect 6328 489960 368572 489988
rect 6328 489948 6334 489960
rect 368566 489948 368572 489960
rect 368624 489948 368630 490000
rect 3418 489880 3424 489932
rect 3476 489920 3482 489932
rect 369854 489920 369860 489932
rect 3476 489892 369860 489920
rect 3476 489880 3482 489892
rect 369854 489880 369860 489892
rect 369912 489880 369918 489932
rect 275922 488452 275928 488504
rect 275980 488492 275986 488504
rect 384114 488492 384120 488504
rect 275980 488464 384120 488492
rect 275980 488452 275986 488464
rect 384114 488452 384120 488464
rect 384172 488452 384178 488504
rect 274542 488384 274548 488436
rect 274600 488424 274606 488436
rect 383194 488424 383200 488436
rect 274600 488396 383200 488424
rect 274600 488384 274606 488396
rect 383194 488384 383200 488396
rect 383252 488384 383258 488436
rect 277118 488316 277124 488368
rect 277176 488356 277182 488368
rect 386138 488356 386144 488368
rect 277176 488328 386144 488356
rect 277176 488316 277182 488328
rect 386138 488316 386144 488328
rect 386196 488316 386202 488368
rect 268286 488248 268292 488300
rect 268344 488288 268350 488300
rect 385862 488288 385868 488300
rect 268344 488260 385868 488288
rect 268344 488248 268350 488260
rect 385862 488248 385868 488260
rect 385920 488248 385926 488300
rect 255222 488180 255228 488232
rect 255280 488220 255286 488232
rect 383378 488220 383384 488232
rect 255280 488192 383384 488220
rect 255280 488180 255286 488192
rect 383378 488180 383384 488192
rect 383436 488180 383442 488232
rect 247586 488112 247592 488164
rect 247644 488152 247650 488164
rect 383102 488152 383108 488164
rect 247644 488124 383108 488152
rect 247644 488112 247650 488124
rect 383102 488112 383108 488124
rect 383160 488112 383166 488164
rect 248874 488044 248880 488096
rect 248932 488084 248938 488096
rect 384666 488084 384672 488096
rect 248932 488056 384672 488084
rect 248932 488044 248938 488056
rect 384666 488044 384672 488056
rect 384724 488044 384730 488096
rect 243722 487976 243728 488028
rect 243780 488016 243786 488028
rect 383010 488016 383016 488028
rect 243780 487988 383016 488016
rect 243780 487976 243786 487988
rect 383010 487976 383016 487988
rect 383068 487976 383074 488028
rect 245010 487908 245016 487960
rect 245068 487948 245074 487960
rect 384574 487948 384580 487960
rect 245068 487920 384580 487948
rect 245068 487908 245074 487920
rect 384574 487908 384580 487920
rect 384632 487908 384638 487960
rect 239858 487840 239864 487892
rect 239916 487880 239922 487892
rect 382918 487880 382924 487892
rect 239916 487852 382924 487880
rect 239916 487840 239922 487852
rect 382918 487840 382924 487852
rect 382976 487840 382982 487892
rect 235902 487772 235908 487824
rect 235960 487812 235966 487824
rect 393958 487812 393964 487824
rect 235960 487784 393964 487812
rect 235960 487772 235966 487784
rect 393958 487772 393964 487784
rect 394016 487772 394022 487824
rect 269252 487704 269258 487756
rect 269310 487744 269316 487756
rect 580902 487744 580908 487756
rect 269310 487716 580908 487744
rect 269310 487704 269316 487716
rect 580902 487704 580908 487716
rect 580960 487704 580966 487756
rect 250162 487636 250168 487688
rect 250220 487676 250226 487688
rect 580350 487676 580356 487688
rect 250220 487648 580356 487676
rect 250220 487636 250226 487648
rect 580350 487636 580356 487648
rect 580408 487636 580414 487688
rect 4706 487568 4712 487620
rect 4764 487608 4770 487620
rect 344002 487608 344008 487620
rect 4764 487580 344008 487608
rect 4764 487568 4770 487580
rect 344002 487568 344008 487580
rect 344060 487568 344066 487620
rect 345290 487608 345296 487620
rect 345251 487580 345296 487608
rect 345290 487568 345296 487580
rect 345348 487568 345354 487620
rect 371234 487608 371240 487620
rect 354646 487580 371240 487608
rect 4982 487500 4988 487552
rect 5040 487540 5046 487552
rect 354646 487540 354674 487580
rect 371234 487568 371240 487580
rect 371292 487568 371298 487620
rect 355594 487540 355600 487552
rect 5040 487512 354674 487540
rect 355555 487512 355600 487540
rect 5040 487500 5046 487512
rect 355594 487500 355600 487512
rect 355652 487500 355658 487552
rect 359458 487540 359464 487552
rect 359419 487512 359464 487540
rect 359458 487500 359464 487512
rect 359516 487500 359522 487552
rect 363414 487540 363420 487552
rect 363375 487512 363420 487540
rect 363414 487500 363420 487512
rect 363472 487500 363478 487552
rect 367278 487540 367284 487552
rect 367239 487512 367284 487540
rect 367278 487500 367284 487512
rect 367336 487500 367342 487552
rect 376294 487540 376300 487552
rect 369136 487512 376300 487540
rect 7742 487432 7748 487484
rect 7800 487472 7806 487484
rect 369136 487472 369164 487512
rect 376294 487500 376300 487512
rect 376352 487500 376358 487552
rect 7800 487444 369164 487472
rect 7800 487432 7806 487444
rect 4890 487364 4896 487416
rect 4948 487404 4954 487416
rect 375006 487404 375012 487416
rect 4948 487376 375012 487404
rect 4948 487364 4954 487376
rect 375006 487364 375012 487376
rect 375064 487364 375070 487416
rect 7558 487296 7564 487348
rect 7616 487336 7622 487348
rect 380158 487336 380164 487348
rect 7616 487308 380164 487336
rect 7616 487296 7622 487308
rect 380158 487296 380164 487308
rect 380216 487296 380222 487348
rect 7650 487228 7656 487280
rect 7708 487268 7714 487280
rect 381446 487268 381452 487280
rect 7708 487240 381452 487268
rect 7708 487228 7714 487240
rect 381446 487228 381452 487240
rect 381504 487228 381510 487280
rect 4798 487160 4804 487212
rect 4856 487200 4862 487212
rect 378870 487200 378876 487212
rect 4856 487172 378876 487200
rect 4856 487160 4862 487172
rect 378870 487160 378876 487172
rect 378928 487160 378934 487212
rect 270862 487092 270868 487144
rect 270920 487132 270926 487144
rect 384206 487132 384212 487144
rect 270920 487104 384212 487132
rect 270920 487092 270926 487104
rect 384206 487092 384212 487104
rect 384264 487092 384270 487144
rect 241146 487024 241152 487076
rect 241204 487064 241210 487076
rect 257890 487064 257896 487076
rect 241204 487036 248414 487064
rect 257851 487036 257896 487064
rect 241204 487024 241210 487036
rect 246298 486956 246304 487008
rect 246356 486956 246362 487008
rect 246316 486180 246344 486956
rect 248386 486588 248414 487036
rect 257890 487024 257896 487036
rect 257948 487024 257954 487076
rect 259270 487024 259276 487076
rect 259328 487064 259334 487076
rect 259328 487036 263088 487064
rect 259328 487024 259334 487036
rect 251266 486956 251272 487008
rect 251324 486956 251330 487008
rect 252554 486996 252560 487008
rect 252515 486968 252560 486996
rect 252554 486956 252560 486968
rect 252612 486956 252618 487008
rect 253842 486996 253848 487008
rect 253803 486968 253848 486996
rect 253842 486956 253848 486968
rect 253900 486956 253906 487008
rect 256602 486956 256608 487008
rect 256660 486996 256666 487008
rect 256660 486968 258074 486996
rect 256660 486956 256666 486968
rect 251284 486724 251312 486956
rect 258046 486792 258074 486968
rect 260558 486956 260564 487008
rect 260616 486956 260622 487008
rect 261846 486996 261852 487008
rect 261807 486968 261852 486996
rect 261846 486956 261852 486968
rect 261904 486956 261910 487008
rect 260576 486860 260604 486956
rect 263060 486928 263088 487036
rect 263134 487024 263140 487076
rect 263192 487064 263198 487076
rect 263192 487036 265848 487064
rect 263192 487024 263198 487036
rect 264422 486996 264428 487008
rect 264383 486968 264428 486996
rect 264422 486956 264428 486968
rect 264480 486956 264486 487008
rect 265710 486996 265716 487008
rect 265671 486968 265716 486996
rect 265710 486956 265716 486968
rect 265768 486956 265774 487008
rect 265820 486996 265848 487036
rect 266998 487024 267004 487076
rect 267056 487064 267062 487076
rect 384942 487064 384948 487076
rect 267056 487036 384948 487064
rect 267056 487024 267062 487036
rect 384942 487024 384948 487036
rect 385000 487024 385006 487076
rect 383562 486996 383568 487008
rect 265820 486968 383568 486996
rect 383562 486956 383568 486968
rect 383620 486956 383626 487008
rect 383470 486928 383476 486940
rect 263060 486900 383476 486928
rect 383470 486888 383476 486900
rect 383528 486888 383534 486940
rect 385770 486860 385776 486872
rect 260576 486832 385776 486860
rect 385770 486820 385776 486832
rect 385828 486820 385834 486872
rect 384850 486792 384856 486804
rect 258046 486764 384856 486792
rect 384850 486752 384856 486764
rect 384908 486752 384914 486804
rect 383286 486724 383292 486736
rect 251284 486696 383292 486724
rect 383286 486684 383292 486696
rect 383344 486684 383350 486736
rect 252557 486659 252615 486665
rect 252557 486625 252569 486659
rect 252603 486656 252615 486659
rect 384758 486656 384764 486668
rect 252603 486628 384764 486656
rect 252603 486625 252615 486628
rect 252557 486619 252615 486625
rect 384758 486616 384764 486628
rect 384816 486616 384822 486668
rect 384390 486588 384396 486600
rect 248386 486560 384396 486588
rect 384390 486548 384396 486560
rect 384448 486548 384454 486600
rect 265713 486523 265771 486529
rect 265713 486489 265725 486523
rect 265759 486520 265771 486523
rect 580718 486520 580724 486532
rect 265759 486492 580724 486520
rect 265759 486489 265771 486492
rect 265713 486483 265771 486489
rect 580718 486480 580724 486492
rect 580776 486480 580782 486532
rect 264425 486455 264483 486461
rect 264425 486421 264437 486455
rect 264471 486452 264483 486455
rect 580810 486452 580816 486464
rect 264471 486424 580816 486452
rect 264471 486421 264483 486424
rect 264425 486415 264483 486421
rect 580810 486412 580816 486424
rect 580868 486412 580874 486464
rect 261849 486387 261907 486393
rect 261849 486353 261861 486387
rect 261895 486384 261907 486387
rect 580626 486384 580632 486396
rect 261895 486356 580632 486384
rect 261895 486353 261907 486356
rect 261849 486347 261907 486353
rect 580626 486344 580632 486356
rect 580684 486344 580690 486396
rect 257893 486319 257951 486325
rect 257893 486285 257905 486319
rect 257939 486316 257951 486319
rect 580534 486316 580540 486328
rect 257939 486288 580540 486316
rect 257939 486285 257951 486288
rect 257893 486279 257951 486285
rect 580534 486276 580540 486288
rect 580592 486276 580598 486328
rect 253845 486251 253903 486257
rect 253845 486217 253857 486251
rect 253891 486248 253903 486251
rect 580442 486248 580448 486260
rect 253891 486220 580448 486248
rect 253891 486217 253903 486220
rect 253845 486211 253903 486217
rect 580442 486208 580448 486220
rect 580500 486208 580506 486260
rect 580258 486180 580264 486192
rect 246316 486152 580264 486180
rect 580258 486140 580264 486152
rect 580316 486140 580322 486192
rect 6638 486072 6644 486124
rect 6696 486112 6702 486124
rect 345293 486115 345351 486121
rect 345293 486112 345305 486115
rect 6696 486084 345305 486112
rect 6696 486072 6702 486084
rect 345293 486081 345305 486084
rect 345339 486081 345351 486115
rect 345293 486075 345351 486081
rect 5166 486004 5172 486056
rect 5224 486044 5230 486056
rect 355597 486047 355655 486053
rect 355597 486044 355609 486047
rect 5224 486016 355609 486044
rect 5224 486004 5230 486016
rect 355597 486013 355609 486016
rect 355643 486013 355655 486047
rect 355597 486007 355655 486013
rect 5074 485936 5080 485988
rect 5132 485976 5138 485988
rect 359461 485979 359519 485985
rect 359461 485976 359473 485979
rect 5132 485948 359473 485976
rect 5132 485936 5138 485948
rect 359461 485945 359473 485948
rect 359507 485945 359519 485979
rect 359461 485939 359519 485945
rect 3694 485868 3700 485920
rect 3752 485908 3758 485920
rect 363417 485911 363475 485917
rect 363417 485908 363429 485911
rect 3752 485880 363429 485908
rect 3752 485868 3758 485880
rect 363417 485877 363429 485880
rect 363463 485877 363475 485911
rect 363417 485871 363475 485877
rect 3510 485800 3516 485852
rect 3568 485840 3574 485852
rect 367281 485843 367339 485849
rect 367281 485840 367293 485843
rect 3568 485812 367293 485840
rect 3568 485800 3574 485812
rect 367281 485809 367293 485812
rect 367327 485809 367339 485843
rect 367281 485803 367339 485809
rect 384114 485732 384120 485784
rect 384172 485772 384178 485784
rect 580166 485772 580172 485784
rect 384172 485744 580172 485772
rect 384172 485732 384178 485744
rect 580166 485732 580172 485744
rect 580224 485732 580230 485784
rect 2774 475668 2780 475720
rect 2832 475708 2838 475720
rect 4706 475708 4712 475720
rect 2832 475680 4712 475708
rect 2832 475668 2838 475680
rect 4706 475668 4712 475680
rect 4764 475668 4770 475720
rect 386138 471928 386144 471980
rect 386196 471968 386202 471980
rect 580166 471968 580172 471980
rect 386196 471940 580172 471968
rect 386196 471928 386202 471940
rect 580166 471928 580172 471940
rect 580224 471928 580230 471980
rect 3234 462680 3240 462732
rect 3292 462720 3298 462732
rect 7926 462720 7932 462732
rect 3292 462692 7932 462720
rect 3292 462680 3298 462692
rect 7926 462680 7932 462692
rect 7984 462680 7990 462732
rect 383194 458124 383200 458176
rect 383252 458164 383258 458176
rect 580166 458164 580172 458176
rect 383252 458136 580172 458164
rect 383252 458124 383258 458136
rect 580166 458124 580172 458136
rect 580224 458124 580230 458176
rect 3234 449556 3240 449608
rect 3292 449596 3298 449608
rect 6638 449596 6644 449608
rect 3292 449568 6644 449596
rect 3292 449556 3298 449568
rect 6638 449556 6644 449568
rect 6696 449556 6702 449608
rect 386046 431876 386052 431928
rect 386104 431916 386110 431928
rect 580166 431916 580172 431928
rect 386104 431888 580172 431916
rect 386104 431876 386110 431888
rect 580166 431876 580172 431888
rect 580224 431876 580230 431928
rect 2774 423580 2780 423632
rect 2832 423620 2838 423632
rect 5442 423620 5448 423632
rect 2832 423592 5448 423620
rect 2832 423580 2838 423592
rect 5442 423580 5448 423592
rect 5500 423580 5506 423632
rect 385954 419432 385960 419484
rect 386012 419472 386018 419484
rect 580166 419472 580172 419484
rect 386012 419444 580172 419472
rect 386012 419432 386018 419444
rect 580166 419432 580172 419444
rect 580224 419432 580230 419484
rect 384206 405628 384212 405680
rect 384264 405668 384270 405680
rect 580166 405668 580172 405680
rect 384264 405640 580172 405668
rect 384264 405628 384270 405640
rect 580166 405628 580172 405640
rect 580224 405628 580230 405680
rect 2774 397536 2780 397588
rect 2832 397576 2838 397588
rect 5350 397576 5356 397588
rect 2832 397548 5356 397576
rect 2832 397536 2838 397548
rect 5350 397536 5356 397548
rect 5408 397536 5414 397588
rect 385862 379448 385868 379500
rect 385920 379488 385926 379500
rect 579982 379488 579988 379500
rect 385920 379460 579988 379488
rect 385920 379448 385926 379460
rect 579982 379448 579988 379460
rect 580040 379448 580046 379500
rect 2774 371424 2780 371476
rect 2832 371464 2838 371476
rect 5258 371464 5264 371476
rect 2832 371436 5264 371464
rect 2832 371424 2838 371436
rect 5258 371424 5264 371436
rect 5316 371424 5322 371476
rect 384942 353200 384948 353252
rect 385000 353240 385006 353252
rect 580166 353240 580172 353252
rect 385000 353212 580172 353240
rect 385000 353200 385006 353212
rect 580166 353200 580172 353212
rect 580224 353200 580230 353252
rect 251220 337764 251226 337816
rect 251278 337804 251284 337816
rect 251542 337804 251548 337816
rect 251278 337776 251548 337804
rect 251278 337764 251284 337776
rect 251542 337764 251548 337776
rect 251600 337764 251606 337816
rect 265020 337764 265026 337816
rect 265078 337804 265084 337816
rect 265250 337804 265256 337816
rect 265078 337776 265256 337804
rect 265078 337764 265084 337776
rect 265250 337764 265256 337776
rect 265308 337764 265314 337816
rect 251192 336756 251680 336784
rect 75822 336676 75828 336728
rect 75880 336716 75886 336728
rect 251192 336716 251220 336756
rect 75880 336688 251220 336716
rect 251652 336716 251680 336756
rect 284294 336744 284300 336796
rect 284352 336784 284358 336796
rect 284662 336784 284668 336796
rect 284352 336756 284668 336784
rect 284352 336744 284358 336756
rect 284662 336744 284668 336756
rect 284720 336744 284726 336796
rect 293954 336744 293960 336796
rect 294012 336784 294018 336796
rect 294782 336784 294788 336796
rect 294012 336756 294788 336784
rect 294012 336744 294018 336756
rect 294782 336744 294788 336756
rect 294840 336744 294846 336796
rect 337930 336744 337936 336796
rect 337988 336744 337994 336796
rect 376110 336744 376116 336796
rect 376168 336784 376174 336796
rect 382185 336787 382243 336793
rect 382185 336784 382197 336787
rect 376168 336756 382197 336784
rect 376168 336744 376174 336756
rect 382185 336753 382197 336756
rect 382231 336753 382243 336787
rect 382185 336747 382243 336753
rect 253750 336716 253756 336728
rect 251652 336688 253756 336716
rect 75880 336676 75886 336688
rect 253750 336676 253756 336688
rect 253808 336676 253814 336728
rect 258166 336676 258172 336728
rect 258224 336716 258230 336728
rect 258534 336716 258540 336728
rect 258224 336688 258540 336716
rect 258224 336676 258230 336688
rect 258534 336676 258540 336688
rect 258592 336676 258598 336728
rect 278314 336716 278320 336728
rect 265360 336688 278320 336716
rect 68922 336608 68928 336660
rect 68980 336648 68986 336660
rect 252002 336648 252008 336660
rect 68980 336620 252008 336648
rect 68980 336608 68986 336620
rect 252002 336608 252008 336620
rect 252060 336608 252066 336660
rect 265360 336648 265388 336688
rect 278314 336676 278320 336688
rect 278372 336676 278378 336728
rect 281534 336676 281540 336728
rect 281592 336716 281598 336728
rect 281902 336716 281908 336728
rect 281592 336688 281908 336716
rect 281592 336676 281598 336688
rect 281902 336676 281908 336688
rect 281960 336676 281966 336728
rect 282270 336676 282276 336728
rect 282328 336716 282334 336728
rect 305178 336716 305184 336728
rect 282328 336688 305184 336716
rect 282328 336676 282334 336688
rect 305178 336676 305184 336688
rect 305236 336676 305242 336728
rect 313366 336676 313372 336728
rect 313424 336716 313430 336728
rect 313550 336716 313556 336728
rect 313424 336688 313556 336716
rect 313424 336676 313430 336688
rect 313550 336676 313556 336688
rect 313608 336676 313614 336728
rect 317782 336676 317788 336728
rect 317840 336716 317846 336728
rect 320818 336716 320824 336728
rect 317840 336688 320824 336716
rect 317840 336676 317846 336688
rect 320818 336676 320824 336688
rect 320876 336676 320882 336728
rect 321186 336676 321192 336728
rect 321244 336716 321250 336728
rect 321462 336716 321468 336728
rect 321244 336688 321468 336716
rect 321244 336676 321250 336688
rect 321462 336676 321468 336688
rect 321520 336676 321526 336728
rect 322014 336676 322020 336728
rect 322072 336716 322078 336728
rect 322750 336716 322756 336728
rect 322072 336688 322756 336716
rect 322072 336676 322078 336688
rect 322750 336676 322756 336688
rect 322808 336676 322814 336728
rect 323854 336676 323860 336728
rect 323912 336716 323918 336728
rect 324222 336716 324228 336728
rect 323912 336688 324228 336716
rect 323912 336676 323918 336688
rect 324222 336676 324228 336688
rect 324280 336676 324286 336728
rect 325234 336676 325240 336728
rect 325292 336716 325298 336728
rect 325510 336716 325516 336728
rect 325292 336688 325516 336716
rect 325292 336676 325298 336688
rect 325510 336676 325516 336688
rect 325568 336676 325574 336728
rect 327626 336676 327632 336728
rect 327684 336716 327690 336728
rect 328270 336716 328276 336728
rect 327684 336688 328276 336716
rect 327684 336676 327690 336688
rect 328270 336676 328276 336688
rect 328328 336676 328334 336728
rect 329466 336676 329472 336728
rect 329524 336716 329530 336728
rect 329742 336716 329748 336728
rect 329524 336688 329748 336716
rect 329524 336676 329530 336688
rect 329742 336676 329748 336688
rect 329800 336676 329806 336728
rect 330662 336676 330668 336728
rect 330720 336716 330726 336728
rect 330846 336716 330852 336728
rect 330720 336688 330852 336716
rect 330720 336676 330726 336688
rect 330846 336676 330852 336688
rect 330904 336676 330910 336728
rect 331858 336676 331864 336728
rect 331916 336716 331922 336728
rect 332318 336716 332324 336728
rect 331916 336688 332324 336716
rect 331916 336676 331922 336688
rect 332318 336676 332324 336688
rect 332376 336676 332382 336728
rect 334894 336676 334900 336728
rect 334952 336716 334958 336728
rect 335262 336716 335268 336728
rect 334952 336688 335268 336716
rect 334952 336676 334958 336688
rect 335262 336676 335268 336688
rect 335320 336676 335326 336728
rect 337654 336676 337660 336728
rect 337712 336716 337718 336728
rect 337948 336716 337976 336744
rect 337712 336688 337976 336716
rect 337712 336676 337718 336688
rect 338758 336676 338764 336728
rect 338816 336716 338822 336728
rect 339126 336716 339132 336728
rect 338816 336688 339132 336716
rect 338816 336676 338822 336688
rect 339126 336676 339132 336688
rect 339184 336676 339190 336728
rect 339218 336676 339224 336728
rect 339276 336716 339282 336728
rect 339402 336716 339408 336728
rect 339276 336688 339408 336716
rect 339276 336676 339282 336688
rect 339402 336676 339408 336688
rect 339460 336676 339466 336728
rect 340506 336676 340512 336728
rect 340564 336716 340570 336728
rect 340782 336716 340788 336728
rect 340564 336688 340788 336716
rect 340564 336676 340570 336688
rect 340782 336676 340788 336688
rect 340840 336676 340846 336728
rect 341426 336676 341432 336728
rect 341484 336716 341490 336728
rect 342162 336716 342168 336728
rect 341484 336688 342168 336716
rect 341484 336676 341490 336688
rect 342162 336676 342168 336688
rect 342220 336676 342226 336728
rect 342622 336676 342628 336728
rect 342680 336716 342686 336728
rect 343358 336716 343364 336728
rect 342680 336688 343364 336716
rect 342680 336676 342686 336688
rect 343358 336676 343364 336688
rect 343416 336676 343422 336728
rect 405090 336716 405096 336728
rect 343652 336688 405096 336716
rect 258046 336620 265388 336648
rect 62022 336540 62028 336592
rect 62080 336580 62086 336592
rect 250162 336580 250168 336592
rect 62080 336552 250168 336580
rect 62080 336540 62086 336552
rect 250162 336540 250168 336552
rect 250220 336540 250226 336592
rect 53742 336472 53748 336524
rect 53800 336512 53806 336524
rect 248414 336512 248420 336524
rect 53800 336484 248420 336512
rect 53800 336472 53806 336484
rect 248414 336472 248420 336484
rect 248472 336472 248478 336524
rect 258046 336512 258074 336620
rect 267642 336608 267648 336660
rect 267700 336648 267706 336660
rect 302234 336648 302240 336660
rect 267700 336620 302240 336648
rect 267700 336608 267706 336620
rect 302234 336608 302240 336620
rect 302292 336608 302298 336660
rect 318794 336608 318800 336660
rect 318852 336648 318858 336660
rect 322198 336648 322204 336660
rect 318852 336620 322204 336648
rect 318852 336608 318858 336620
rect 322198 336608 322204 336620
rect 322256 336608 322262 336660
rect 324682 336608 324688 336660
rect 324740 336648 324746 336660
rect 325326 336648 325332 336660
rect 324740 336620 325332 336648
rect 324740 336608 324746 336620
rect 325326 336608 325332 336620
rect 325384 336608 325390 336660
rect 326430 336608 326436 336660
rect 326488 336648 326494 336660
rect 326798 336648 326804 336660
rect 326488 336620 326804 336648
rect 326488 336608 326494 336620
rect 326798 336608 326804 336620
rect 326856 336608 326862 336660
rect 328822 336608 328828 336660
rect 328880 336648 328886 336660
rect 329650 336648 329656 336660
rect 328880 336620 329656 336648
rect 328880 336608 328886 336620
rect 329650 336608 329656 336620
rect 329708 336608 329714 336660
rect 330018 336608 330024 336660
rect 330076 336648 330082 336660
rect 330938 336648 330944 336660
rect 330076 336620 330944 336648
rect 330076 336608 330082 336620
rect 330938 336608 330944 336620
rect 330996 336608 331002 336660
rect 331950 336608 331956 336660
rect 332008 336648 332014 336660
rect 332502 336648 332508 336660
rect 332008 336620 332508 336648
rect 332008 336608 332014 336620
rect 332502 336608 332508 336620
rect 332560 336608 332566 336660
rect 334250 336608 334256 336660
rect 334308 336648 334314 336660
rect 335078 336648 335084 336660
rect 334308 336620 335084 336648
rect 334308 336608 334314 336620
rect 335078 336608 335084 336620
rect 335136 336608 335142 336660
rect 339954 336608 339960 336660
rect 340012 336648 340018 336660
rect 340690 336648 340696 336660
rect 340012 336620 340696 336648
rect 340012 336608 340018 336620
rect 340690 336608 340696 336620
rect 340748 336608 340754 336660
rect 342898 336608 342904 336660
rect 342956 336648 342962 336660
rect 343542 336648 343548 336660
rect 342956 336620 343548 336648
rect 342956 336608 342962 336620
rect 343542 336608 343548 336620
rect 343600 336608 343606 336660
rect 263502 336540 263508 336592
rect 263560 336580 263566 336592
rect 301314 336580 301320 336592
rect 263560 336552 301320 336580
rect 263560 336540 263566 336552
rect 301314 336540 301320 336552
rect 301372 336540 301378 336592
rect 311158 336540 311164 336592
rect 311216 336580 311222 336592
rect 311894 336580 311900 336592
rect 311216 336552 311900 336580
rect 311216 336540 311222 336552
rect 311894 336540 311900 336552
rect 311952 336540 311958 336592
rect 318058 336540 318064 336592
rect 318116 336580 318122 336592
rect 318610 336580 318616 336592
rect 318116 336552 318616 336580
rect 318116 336540 318122 336552
rect 318610 336540 318616 336552
rect 318668 336540 318674 336592
rect 324958 336540 324964 336592
rect 325016 336580 325022 336592
rect 325602 336580 325608 336592
rect 325016 336552 325608 336580
rect 325016 336540 325022 336552
rect 325602 336540 325608 336552
rect 325660 336540 325666 336592
rect 325878 336540 325884 336592
rect 325936 336580 325942 336592
rect 326982 336580 326988 336592
rect 325936 336552 326988 336580
rect 325936 336540 325942 336552
rect 326982 336540 326988 336552
rect 327040 336540 327046 336592
rect 337562 336540 337568 336592
rect 337620 336580 337626 336592
rect 338758 336580 338764 336592
rect 337620 336552 338764 336580
rect 337620 336540 337626 336552
rect 338758 336540 338764 336552
rect 338816 336540 338822 336592
rect 341150 336540 341156 336592
rect 341208 336580 341214 336592
rect 343652 336580 343680 336688
rect 405090 336676 405096 336688
rect 405148 336676 405154 336728
rect 343818 336608 343824 336660
rect 343876 336648 343882 336660
rect 344922 336648 344928 336660
rect 343876 336620 344928 336648
rect 343876 336608 343882 336620
rect 344922 336608 344928 336620
rect 344980 336608 344986 336660
rect 345290 336608 345296 336660
rect 345348 336648 345354 336660
rect 346026 336648 346032 336660
rect 345348 336620 346032 336648
rect 345348 336608 345354 336620
rect 346026 336608 346032 336620
rect 346084 336608 346090 336660
rect 346854 336608 346860 336660
rect 346912 336648 346918 336660
rect 347498 336648 347504 336660
rect 346912 336620 347504 336648
rect 346912 336608 346918 336620
rect 347498 336608 347504 336620
rect 347556 336608 347562 336660
rect 348602 336608 348608 336660
rect 348660 336648 348666 336660
rect 349062 336648 349068 336660
rect 348660 336620 349068 336648
rect 348660 336608 348666 336620
rect 349062 336608 349068 336620
rect 349120 336608 349126 336660
rect 349798 336608 349804 336660
rect 349856 336648 349862 336660
rect 350258 336648 350264 336660
rect 349856 336620 350264 336648
rect 349856 336608 349862 336620
rect 350258 336608 350264 336620
rect 350316 336608 350322 336660
rect 351270 336608 351276 336660
rect 351328 336648 351334 336660
rect 351730 336648 351736 336660
rect 351328 336620 351736 336648
rect 351328 336608 351334 336620
rect 351730 336608 351736 336620
rect 351788 336608 351794 336660
rect 352926 336608 352932 336660
rect 352984 336648 352990 336660
rect 353110 336648 353116 336660
rect 352984 336620 353116 336648
rect 352984 336608 352990 336620
rect 353110 336608 353116 336620
rect 353168 336608 353174 336660
rect 354030 336608 354036 336660
rect 354088 336648 354094 336660
rect 354490 336648 354496 336660
rect 354088 336620 354496 336648
rect 354088 336608 354094 336620
rect 354490 336608 354496 336620
rect 354548 336608 354554 336660
rect 417418 336648 417424 336660
rect 354646 336620 417424 336648
rect 341208 336552 343680 336580
rect 341208 336540 341214 336552
rect 345934 336540 345940 336592
rect 345992 336580 345998 336592
rect 346210 336580 346216 336592
rect 345992 336552 346216 336580
rect 345992 336540 345998 336552
rect 346210 336540 346216 336552
rect 346268 336540 346274 336592
rect 347406 336540 347412 336592
rect 347464 336580 347470 336592
rect 347682 336580 347688 336592
rect 347464 336552 347688 336580
rect 347464 336540 347470 336552
rect 347682 336540 347688 336552
rect 347740 336540 347746 336592
rect 348050 336540 348056 336592
rect 348108 336580 348114 336592
rect 348878 336580 348884 336592
rect 348108 336552 348884 336580
rect 348108 336540 348114 336552
rect 348878 336540 348884 336552
rect 348936 336540 348942 336592
rect 349522 336540 349528 336592
rect 349580 336580 349586 336592
rect 350442 336580 350448 336592
rect 349580 336552 350448 336580
rect 349580 336540 349586 336552
rect 350442 336540 350448 336552
rect 350500 336540 350506 336592
rect 350718 336540 350724 336592
rect 350776 336580 350782 336592
rect 351546 336580 351552 336592
rect 350776 336552 351552 336580
rect 350776 336540 350782 336552
rect 351546 336540 351552 336552
rect 351604 336540 351610 336592
rect 351917 336583 351975 336589
rect 351917 336549 351929 336583
rect 351963 336580 351975 336583
rect 354646 336580 354674 336620
rect 417418 336608 417424 336620
rect 417476 336608 417482 336660
rect 351963 336552 354674 336580
rect 351963 336549 351975 336552
rect 351917 336543 351975 336549
rect 354858 336540 354864 336592
rect 354916 336580 354922 336592
rect 355686 336580 355692 336592
rect 354916 336552 355692 336580
rect 354916 336540 354922 336552
rect 355686 336540 355692 336552
rect 355744 336540 355750 336592
rect 359642 336540 359648 336592
rect 359700 336580 359706 336592
rect 360102 336580 360108 336592
rect 359700 336552 360108 336580
rect 359700 336540 359706 336552
rect 360102 336540 360108 336552
rect 360160 336540 360166 336592
rect 360562 336540 360568 336592
rect 360620 336580 360626 336592
rect 361298 336580 361304 336592
rect 360620 336552 361304 336580
rect 360620 336540 360626 336552
rect 361298 336540 361304 336552
rect 361356 336540 361362 336592
rect 362402 336540 362408 336592
rect 362460 336580 362466 336592
rect 362678 336580 362684 336592
rect 362460 336552 362684 336580
rect 362460 336540 362466 336552
rect 362678 336540 362684 336552
rect 362736 336540 362742 336592
rect 363230 336540 363236 336592
rect 363288 336580 363294 336592
rect 364150 336580 364156 336592
rect 363288 336552 364156 336580
rect 363288 336540 363294 336552
rect 364150 336540 364156 336552
rect 364208 336540 364214 336592
rect 364245 336583 364303 336589
rect 364245 336549 364257 336583
rect 364291 336580 364303 336583
rect 425698 336580 425704 336592
rect 364291 336552 425704 336580
rect 364291 336549 364303 336552
rect 364245 336543 364303 336549
rect 425698 336540 425704 336552
rect 425756 336540 425762 336592
rect 253216 336484 258074 336512
rect 265437 336515 265495 336521
rect 42702 336404 42708 336456
rect 42760 336444 42766 336456
rect 245378 336444 245384 336456
rect 42760 336416 245384 336444
rect 42760 336404 42766 336416
rect 245378 336404 245384 336416
rect 245436 336404 245442 336456
rect 37182 336336 37188 336388
rect 37240 336376 37246 336388
rect 243906 336376 243912 336388
rect 37240 336348 243912 336376
rect 37240 336336 37246 336348
rect 243906 336336 243912 336348
rect 243964 336336 243970 336388
rect 245010 336336 245016 336388
rect 245068 336376 245074 336388
rect 253216 336376 253244 336484
rect 265437 336481 265449 336515
rect 265483 336512 265495 336515
rect 300394 336512 300400 336524
rect 265483 336484 300400 336512
rect 265483 336481 265495 336484
rect 265437 336475 265495 336481
rect 300394 336472 300400 336484
rect 300452 336472 300458 336524
rect 307662 336472 307668 336524
rect 307720 336512 307726 336524
rect 312354 336512 312360 336524
rect 307720 336484 312360 336512
rect 307720 336472 307726 336484
rect 312354 336472 312360 336484
rect 312412 336472 312418 336524
rect 316586 336472 316592 336524
rect 316644 336512 316650 336524
rect 320910 336512 320916 336524
rect 316644 336484 320916 336512
rect 316644 336472 316650 336484
rect 320910 336472 320916 336484
rect 320968 336472 320974 336524
rect 341978 336472 341984 336524
rect 342036 336512 342042 336524
rect 416038 336512 416044 336524
rect 342036 336484 416044 336512
rect 342036 336472 342042 336484
rect 416038 336472 416044 336484
rect 416096 336472 416102 336524
rect 254578 336404 254584 336456
rect 254636 336444 254642 336456
rect 296806 336444 296812 336456
rect 254636 336416 296812 336444
rect 254636 336404 254642 336416
rect 296806 336404 296812 336416
rect 296864 336404 296870 336456
rect 316862 336404 316868 336456
rect 316920 336444 316926 336456
rect 322382 336444 322388 336456
rect 316920 336416 322388 336444
rect 316920 336404 316926 336416
rect 322382 336404 322388 336416
rect 322440 336404 322446 336456
rect 344738 336404 344744 336456
rect 344796 336444 344802 336456
rect 429838 336444 429844 336456
rect 344796 336416 429844 336444
rect 344796 336404 344802 336416
rect 429838 336404 429844 336416
rect 429896 336404 429902 336456
rect 245068 336348 253244 336376
rect 245068 336336 245074 336348
rect 256602 336336 256608 336388
rect 256660 336376 256666 336388
rect 299566 336376 299572 336388
rect 256660 336348 299572 336376
rect 256660 336336 256666 336348
rect 299566 336336 299572 336348
rect 299624 336336 299630 336388
rect 319990 336336 319996 336388
rect 320048 336376 320054 336388
rect 335722 336376 335728 336388
rect 320048 336348 335728 336376
rect 320048 336336 320054 336348
rect 335722 336336 335728 336348
rect 335780 336336 335786 336388
rect 345658 336336 345664 336388
rect 345716 336376 345722 336388
rect 346302 336376 346308 336388
rect 345716 336348 346308 336376
rect 345716 336336 345722 336348
rect 346302 336336 346308 336348
rect 346360 336336 346366 336388
rect 350994 336336 351000 336388
rect 351052 336376 351058 336388
rect 351822 336376 351828 336388
rect 351052 336348 351828 336376
rect 351052 336336 351058 336348
rect 351822 336336 351828 336348
rect 351880 336336 351886 336388
rect 352009 336379 352067 336385
rect 352009 336345 352021 336379
rect 352055 336376 352067 336379
rect 432598 336376 432604 336388
rect 352055 336348 432604 336376
rect 352055 336345 352067 336348
rect 352009 336339 352067 336345
rect 432598 336336 432604 336348
rect 432656 336336 432662 336388
rect 44082 336268 44088 336320
rect 44140 336308 44146 336320
rect 245654 336308 245660 336320
rect 44140 336280 245660 336308
rect 44140 336268 44146 336280
rect 245654 336268 245660 336280
rect 245712 336268 245718 336320
rect 246390 336268 246396 336320
rect 246448 336308 246454 336320
rect 290274 336308 290280 336320
rect 246448 336280 290280 336308
rect 246448 336268 246454 336280
rect 290274 336268 290280 336280
rect 290332 336268 290338 336320
rect 315390 336268 315396 336320
rect 315448 336308 315454 336320
rect 316310 336308 316316 336320
rect 315448 336280 316316 336308
rect 315448 336268 315454 336280
rect 316310 336268 316316 336280
rect 316368 336268 316374 336320
rect 319898 336268 319904 336320
rect 319956 336308 319962 336320
rect 334434 336308 334440 336320
rect 319956 336280 334440 336308
rect 319956 336268 319962 336280
rect 334434 336268 334440 336280
rect 334492 336268 334498 336320
rect 344094 336268 344100 336320
rect 344152 336308 344158 336320
rect 344738 336308 344744 336320
rect 344152 336280 344744 336308
rect 344152 336268 344158 336280
rect 344738 336268 344744 336280
rect 344796 336268 344802 336320
rect 349154 336268 349160 336320
rect 349212 336308 349218 336320
rect 351917 336311 351975 336317
rect 351917 336308 351929 336311
rect 349212 336280 351929 336308
rect 349212 336268 349218 336280
rect 351917 336277 351929 336280
rect 351963 336277 351975 336311
rect 351917 336271 351975 336277
rect 352834 336268 352840 336320
rect 352892 336308 352898 336320
rect 353202 336308 353208 336320
rect 352892 336280 353208 336308
rect 352892 336268 352898 336280
rect 353202 336268 353208 336280
rect 353260 336268 353266 336320
rect 353297 336311 353355 336317
rect 353297 336277 353309 336311
rect 353343 336308 353355 336311
rect 436738 336308 436744 336320
rect 353343 336280 436744 336308
rect 353343 336277 353355 336280
rect 353297 336271 353355 336277
rect 436738 336268 436744 336280
rect 436796 336268 436802 336320
rect 35802 336200 35808 336252
rect 35860 336240 35866 336252
rect 243630 336240 243636 336252
rect 35860 336212 243636 336240
rect 35860 336200 35866 336212
rect 243630 336200 243636 336212
rect 243688 336200 243694 336252
rect 251818 336200 251824 336252
rect 251876 336240 251882 336252
rect 295978 336240 295984 336252
rect 251876 336212 295984 336240
rect 251876 336200 251882 336212
rect 295978 336200 295984 336212
rect 296036 336200 296042 336252
rect 319254 336200 319260 336252
rect 319312 336240 319318 336252
rect 324958 336240 324964 336252
rect 319312 336212 324964 336240
rect 319312 336200 319318 336212
rect 324958 336200 324964 336212
rect 325016 336200 325022 336252
rect 350074 336200 350080 336252
rect 350132 336240 350138 336252
rect 440878 336240 440884 336252
rect 350132 336212 440884 336240
rect 350132 336200 350138 336212
rect 440878 336200 440884 336212
rect 440936 336200 440942 336252
rect 28902 336132 28908 336184
rect 28960 336172 28966 336184
rect 241790 336172 241796 336184
rect 28960 336144 241796 336172
rect 28960 336132 28966 336144
rect 241790 336132 241796 336144
rect 241848 336132 241854 336184
rect 244918 336132 244924 336184
rect 244976 336172 244982 336184
rect 290090 336172 290096 336184
rect 244976 336144 290096 336172
rect 244976 336132 244982 336144
rect 290090 336132 290096 336144
rect 290148 336132 290154 336184
rect 320726 336132 320732 336184
rect 320784 336172 320790 336184
rect 338574 336172 338580 336184
rect 320784 336144 338580 336172
rect 320784 336132 320790 336144
rect 338574 336132 338580 336144
rect 338632 336132 338638 336184
rect 346394 336132 346400 336184
rect 346452 336172 346458 336184
rect 351825 336175 351883 336181
rect 351825 336172 351837 336175
rect 346452 336144 351837 336172
rect 346452 336132 346458 336144
rect 351825 336141 351837 336144
rect 351871 336141 351883 336175
rect 351825 336135 351883 336141
rect 351914 336132 351920 336184
rect 351972 336172 351978 336184
rect 443638 336172 443644 336184
rect 351972 336144 443644 336172
rect 351972 336132 351978 336144
rect 443638 336132 443644 336144
rect 443696 336132 443702 336184
rect 19242 336064 19248 336116
rect 19300 336104 19306 336116
rect 239398 336104 239404 336116
rect 19300 336076 239404 336104
rect 19300 336064 19306 336076
rect 239398 336064 239404 336076
rect 239456 336064 239462 336116
rect 252462 336064 252468 336116
rect 252520 336104 252526 336116
rect 298646 336104 298652 336116
rect 252520 336076 298652 336104
rect 252520 336064 252526 336076
rect 298646 336064 298652 336076
rect 298704 336064 298710 336116
rect 315942 336064 315948 336116
rect 316000 336104 316006 336116
rect 318886 336104 318892 336116
rect 316000 336076 318892 336104
rect 316000 336064 316006 336076
rect 318886 336064 318892 336076
rect 318944 336064 318950 336116
rect 321094 336064 321100 336116
rect 321152 336104 321158 336116
rect 339862 336104 339868 336116
rect 321152 336076 339868 336104
rect 321152 336064 321158 336076
rect 339862 336064 339868 336076
rect 339920 336064 339926 336116
rect 348326 336064 348332 336116
rect 348384 336104 348390 336116
rect 353297 336107 353355 336113
rect 353297 336104 353309 336107
rect 348384 336076 353309 336104
rect 348384 336064 348390 336076
rect 353297 336073 353309 336076
rect 353343 336073 353355 336107
rect 353297 336067 353355 336073
rect 353662 336064 353668 336116
rect 353720 336104 353726 336116
rect 447778 336104 447784 336116
rect 353720 336076 447784 336104
rect 353720 336064 353726 336076
rect 447778 336064 447784 336076
rect 447836 336064 447842 336116
rect 20622 335996 20628 336048
rect 20680 336036 20686 336048
rect 240134 336036 240140 336048
rect 20680 336008 240140 336036
rect 20680 335996 20686 336008
rect 240134 335996 240140 336008
rect 240192 335996 240198 336048
rect 249058 335996 249064 336048
rect 249116 336036 249122 336048
rect 296530 336036 296536 336048
rect 249116 336008 296536 336036
rect 249116 335996 249122 336008
rect 296530 335996 296536 336008
rect 296588 335996 296594 336048
rect 303522 335996 303528 336048
rect 303580 336036 303586 336048
rect 311526 336036 311532 336048
rect 303580 336008 311532 336036
rect 303580 335996 303586 336008
rect 311526 335996 311532 336008
rect 311584 335996 311590 336048
rect 316126 335996 316132 336048
rect 316184 336036 316190 336048
rect 317966 336036 317972 336048
rect 316184 336008 317972 336036
rect 316184 335996 316190 336008
rect 317966 335996 317972 336008
rect 318024 335996 318030 336048
rect 322842 335996 322848 336048
rect 322900 336036 322906 336048
rect 346762 336036 346768 336048
rect 322900 336008 346768 336036
rect 322900 335996 322906 336008
rect 346762 335996 346768 336008
rect 346820 335996 346826 336048
rect 357894 335996 357900 336048
rect 357952 336036 357958 336048
rect 358722 336036 358728 336048
rect 357952 336008 358728 336036
rect 357952 335996 357958 336008
rect 358722 335996 358728 336008
rect 358780 335996 358786 336048
rect 359090 335996 359096 336048
rect 359148 336036 359154 336048
rect 359918 336036 359924 336048
rect 359148 336008 359924 336036
rect 359148 335996 359154 336008
rect 359918 335996 359924 336008
rect 359976 335996 359982 336048
rect 361758 335996 361764 336048
rect 361816 336036 361822 336048
rect 362586 336036 362592 336048
rect 361816 336008 362592 336036
rect 361816 335996 361822 336008
rect 362586 335996 362592 336008
rect 362644 335996 362650 336048
rect 362681 336039 362739 336045
rect 362681 336005 362693 336039
rect 362727 336036 362739 336039
rect 450538 336036 450544 336048
rect 362727 336008 450544 336036
rect 362727 336005 362739 336008
rect 362681 335999 362739 336005
rect 450538 335996 450544 336008
rect 450596 335996 450602 336048
rect 82722 335928 82728 335980
rect 82780 335968 82786 335980
rect 255590 335968 255596 335980
rect 82780 335940 255596 335968
rect 82780 335928 82786 335940
rect 255590 335928 255596 335940
rect 255648 335928 255654 335980
rect 260742 335928 260748 335980
rect 260800 335968 260806 335980
rect 265437 335971 265495 335977
rect 265437 335968 265449 335971
rect 260800 335940 265449 335968
rect 260800 335928 260806 335940
rect 265437 335937 265449 335940
rect 265483 335937 265495 335971
rect 265437 335931 265495 335937
rect 269022 335928 269028 335980
rect 269080 335968 269086 335980
rect 302786 335968 302792 335980
rect 269080 335940 302792 335968
rect 269080 335928 269086 335940
rect 302786 335928 302792 335940
rect 302844 335928 302850 335980
rect 323210 335928 323216 335980
rect 323268 335968 323274 335980
rect 324130 335968 324136 335980
rect 323268 335940 324136 335968
rect 323268 335928 323274 335940
rect 324130 335928 324136 335940
rect 324188 335928 324194 335980
rect 337286 335928 337292 335980
rect 337344 335968 337350 335980
rect 337746 335968 337752 335980
rect 337344 335940 337752 335968
rect 337344 335928 337350 335940
rect 337746 335928 337752 335940
rect 337804 335928 337810 335980
rect 343174 335928 343180 335980
rect 343232 335968 343238 335980
rect 343450 335968 343456 335980
rect 343232 335940 343456 335968
rect 343232 335928 343238 335940
rect 343450 335928 343456 335940
rect 343508 335928 343514 335980
rect 391198 335968 391204 335980
rect 343560 335940 391204 335968
rect 93762 335860 93768 335912
rect 93820 335900 93826 335912
rect 258350 335900 258356 335912
rect 93820 335872 258356 335900
rect 93820 335860 93826 335872
rect 258350 335860 258356 335872
rect 258408 335860 258414 335912
rect 271230 335860 271236 335912
rect 271288 335900 271294 335912
rect 301958 335900 301964 335912
rect 271288 335872 301964 335900
rect 271288 335860 271294 335872
rect 301958 335860 301964 335872
rect 302016 335860 302022 335912
rect 340230 335860 340236 335912
rect 340288 335900 340294 335912
rect 343560 335900 343588 335940
rect 391198 335928 391204 335940
rect 391256 335928 391262 335980
rect 340288 335872 343588 335900
rect 344986 335872 379560 335900
rect 340288 335860 340294 335872
rect 86862 335792 86868 335844
rect 86920 335832 86926 335844
rect 256418 335832 256424 335844
rect 86920 335804 256424 335832
rect 86920 335792 86926 335804
rect 256418 335792 256424 335804
rect 256476 335792 256482 335844
rect 274542 335792 274548 335844
rect 274600 335832 274606 335844
rect 303982 335832 303988 335844
rect 274600 335804 303988 335832
rect 274600 335792 274606 335804
rect 303982 335792 303988 335804
rect 304040 335792 304046 335844
rect 327350 335792 327356 335844
rect 327408 335832 327414 335844
rect 328086 335832 328092 335844
rect 327408 335804 328092 335832
rect 327408 335792 327414 335804
rect 328086 335792 328092 335804
rect 328144 335792 328150 335844
rect 333054 335792 333060 335844
rect 333112 335832 333118 335844
rect 333882 335832 333888 335844
rect 333112 335804 333888 335832
rect 333112 335792 333118 335804
rect 333882 335792 333888 335804
rect 333940 335792 333946 335844
rect 338482 335792 338488 335844
rect 338540 335832 338546 335844
rect 344986 335832 345014 335872
rect 338540 335804 345014 335832
rect 338540 335792 338546 335804
rect 362034 335792 362040 335844
rect 362092 335832 362098 335844
rect 362862 335832 362868 335844
rect 362092 335804 362868 335832
rect 362092 335792 362098 335804
rect 362862 335792 362868 335804
rect 362920 335792 362926 335844
rect 364242 335792 364248 335844
rect 364300 335832 364306 335844
rect 364300 335792 364334 335832
rect 366266 335792 366272 335844
rect 366324 335832 366330 335844
rect 366726 335832 366732 335844
rect 366324 335804 366732 335832
rect 366324 335792 366330 335804
rect 366726 335792 366732 335804
rect 366784 335792 366790 335844
rect 366910 335792 366916 335844
rect 366968 335832 366974 335844
rect 366968 335804 367416 335832
rect 366968 335792 366974 335804
rect 100662 335724 100668 335776
rect 100720 335764 100726 335776
rect 260006 335764 260012 335776
rect 100720 335736 260012 335764
rect 100720 335724 100726 335736
rect 260006 335724 260012 335736
rect 260064 335724 260070 335776
rect 285582 335724 285588 335776
rect 285640 335764 285646 335776
rect 306742 335764 306748 335776
rect 285640 335736 306748 335764
rect 285640 335724 285646 335736
rect 306742 335724 306748 335736
rect 306800 335724 306806 335776
rect 335538 335724 335544 335776
rect 335596 335764 335602 335776
rect 336550 335764 336556 335776
rect 335596 335736 336556 335764
rect 335596 335724 335602 335736
rect 336550 335724 336556 335736
rect 336608 335724 336614 335776
rect 356422 335724 356428 335776
rect 356480 335764 356486 335776
rect 364153 335767 364211 335773
rect 364153 335764 364165 335767
rect 356480 335736 364165 335764
rect 356480 335724 356486 335736
rect 364153 335733 364165 335736
rect 364199 335733 364211 335767
rect 364153 335727 364211 335733
rect 107562 335656 107568 335708
rect 107620 335696 107626 335708
rect 261846 335696 261852 335708
rect 107620 335668 261852 335696
rect 107620 335656 107626 335668
rect 261846 335656 261852 335668
rect 261904 335656 261910 335708
rect 288342 335656 288348 335708
rect 288400 335696 288406 335708
rect 307754 335696 307760 335708
rect 288400 335668 307760 335696
rect 288400 335656 288406 335668
rect 307754 335656 307760 335668
rect 307812 335656 307818 335708
rect 330386 335656 330392 335708
rect 330444 335696 330450 335708
rect 331122 335696 331128 335708
rect 330444 335668 331128 335696
rect 330444 335656 330450 335668
rect 331122 335656 331128 335668
rect 331180 335656 331186 335708
rect 331582 335656 331588 335708
rect 331640 335696 331646 335708
rect 332226 335696 332232 335708
rect 331640 335668 332232 335696
rect 331640 335656 331646 335668
rect 332226 335656 332232 335668
rect 332284 335656 332290 335708
rect 336918 335656 336924 335708
rect 336976 335696 336982 335708
rect 337930 335696 337936 335708
rect 336976 335668 337936 335696
rect 336976 335656 336982 335668
rect 337930 335656 337936 335668
rect 337988 335656 337994 335708
rect 355226 335656 355232 335708
rect 355284 335696 355290 335708
rect 355870 335696 355876 335708
rect 355284 335668 355876 335696
rect 355284 335656 355290 335668
rect 355870 335656 355876 335668
rect 355928 335656 355934 335708
rect 361206 335656 361212 335708
rect 361264 335696 361270 335708
rect 361482 335696 361488 335708
rect 361264 335668 361488 335696
rect 361264 335656 361270 335668
rect 361482 335656 361488 335668
rect 361540 335656 361546 335708
rect 114462 335588 114468 335640
rect 114520 335628 114526 335640
rect 263594 335628 263600 335640
rect 114520 335600 263600 335628
rect 114520 335588 114526 335600
rect 263594 335588 263600 335600
rect 263652 335588 263658 335640
rect 286962 335588 286968 335640
rect 287020 335628 287026 335640
rect 307294 335628 307300 335640
rect 287020 335600 307300 335628
rect 287020 335588 287026 335600
rect 307294 335588 307300 335600
rect 307352 335588 307358 335640
rect 315114 335588 315120 335640
rect 315172 335628 315178 335640
rect 316126 335628 316132 335640
rect 315172 335600 316132 335628
rect 315172 335588 315178 335600
rect 316126 335588 316132 335600
rect 316184 335588 316190 335640
rect 355502 335588 355508 335640
rect 355560 335628 355566 335640
rect 362681 335631 362739 335637
rect 362681 335628 362693 335631
rect 355560 335600 362693 335628
rect 355560 335588 355566 335600
rect 362681 335597 362693 335600
rect 362727 335597 362739 335631
rect 362681 335591 362739 335597
rect 121362 335520 121368 335572
rect 121420 335560 121426 335572
rect 265434 335560 265440 335572
rect 121420 335532 265440 335560
rect 121420 335520 121426 335532
rect 265434 335520 265440 335532
rect 265492 335520 265498 335572
rect 289722 335520 289728 335572
rect 289780 335560 289786 335572
rect 307938 335560 307944 335572
rect 289780 335532 307944 335560
rect 289780 335520 289786 335532
rect 307938 335520 307944 335532
rect 307996 335520 308002 335572
rect 319622 335520 319628 335572
rect 319680 335560 319686 335572
rect 320082 335560 320088 335572
rect 319680 335532 320088 335560
rect 319680 335520 319686 335532
rect 320082 335520 320088 335532
rect 320140 335520 320146 335572
rect 364306 335560 364334 335792
rect 366542 335724 366548 335776
rect 366600 335764 366606 335776
rect 367002 335764 367008 335776
rect 366600 335736 367008 335764
rect 366600 335724 366606 335736
rect 367002 335724 367008 335736
rect 367060 335724 367066 335776
rect 365990 335656 365996 335708
rect 366048 335696 366054 335708
rect 366910 335696 366916 335708
rect 366048 335668 366916 335696
rect 366048 335656 366054 335668
rect 366910 335656 366916 335668
rect 366968 335656 366974 335708
rect 367388 335696 367416 335804
rect 367738 335792 367744 335844
rect 367796 335832 367802 335844
rect 368198 335832 368204 335844
rect 367796 335804 368204 335832
rect 367796 335792 367802 335804
rect 368198 335792 368204 335804
rect 368256 335792 368262 335844
rect 369210 335792 369216 335844
rect 369268 335832 369274 335844
rect 369670 335832 369676 335844
rect 369268 335804 369676 335832
rect 369268 335792 369274 335804
rect 369670 335792 369676 335804
rect 369728 335792 369734 335844
rect 370774 335792 370780 335844
rect 370832 335832 370838 335844
rect 370832 335804 379468 335832
rect 370832 335792 370838 335804
rect 367462 335724 367468 335776
rect 367520 335764 367526 335776
rect 368290 335764 368296 335776
rect 367520 335736 368296 335764
rect 367520 335724 367526 335736
rect 368290 335724 368296 335736
rect 368348 335724 368354 335776
rect 368658 335724 368664 335776
rect 368716 335764 368722 335776
rect 369486 335764 369492 335776
rect 368716 335736 369492 335764
rect 368716 335724 368722 335736
rect 369486 335724 369492 335736
rect 369544 335724 369550 335776
rect 372522 335724 372528 335776
rect 372580 335764 372586 335776
rect 377493 335767 377551 335773
rect 377493 335764 377505 335767
rect 372580 335736 377505 335764
rect 372580 335724 372586 335736
rect 377493 335733 377505 335736
rect 377539 335733 377551 335767
rect 377493 335727 377551 335733
rect 378778 335724 378784 335776
rect 378836 335764 378842 335776
rect 379238 335764 379244 335776
rect 378836 335736 379244 335764
rect 378836 335724 378842 335736
rect 379238 335724 379244 335736
rect 379296 335724 379302 335776
rect 379333 335699 379391 335705
rect 379333 335696 379345 335699
rect 367388 335668 379345 335696
rect 379333 335665 379345 335668
rect 379379 335665 379391 335699
rect 379440 335696 379468 335804
rect 379532 335764 379560 335872
rect 380342 335860 380348 335912
rect 380400 335900 380406 335912
rect 380618 335900 380624 335912
rect 380400 335872 380624 335900
rect 380400 335860 380406 335872
rect 380618 335860 380624 335872
rect 380676 335860 380682 335912
rect 380713 335903 380771 335909
rect 380713 335869 380725 335903
rect 380759 335900 380771 335903
rect 380759 335872 380940 335900
rect 380759 335869 380771 335872
rect 380713 335863 380771 335869
rect 379974 335792 379980 335844
rect 380032 335832 380038 335844
rect 380802 335832 380808 335844
rect 380032 335804 380808 335832
rect 380032 335792 380038 335804
rect 380802 335792 380808 335804
rect 380860 335792 380866 335844
rect 380912 335832 380940 335872
rect 381170 335860 381176 335912
rect 381228 335900 381234 335912
rect 382090 335900 382096 335912
rect 381228 335872 382096 335900
rect 381228 335860 381234 335872
rect 382090 335860 382096 335872
rect 382148 335860 382154 335912
rect 382185 335903 382243 335909
rect 382185 335869 382197 335903
rect 382231 335900 382243 335903
rect 382231 335872 383654 335900
rect 382231 335869 382243 335872
rect 382185 335863 382243 335869
rect 383194 335832 383200 335844
rect 380912 335804 383200 335832
rect 383194 335792 383200 335804
rect 383252 335792 383258 335844
rect 383626 335832 383654 335872
rect 411898 335832 411904 335844
rect 383626 335804 411904 335832
rect 411898 335792 411904 335804
rect 411956 335792 411962 335844
rect 380621 335767 380679 335773
rect 380621 335764 380633 335767
rect 379532 335736 380633 335764
rect 380621 335733 380633 335736
rect 380667 335733 380679 335767
rect 380621 335727 380679 335733
rect 380713 335767 380771 335773
rect 380713 335733 380725 335767
rect 380759 335764 380771 335767
rect 413278 335764 413284 335776
rect 380759 335736 413284 335764
rect 380759 335733 380771 335736
rect 380713 335727 380771 335733
rect 413278 335724 413284 335736
rect 413336 335724 413342 335776
rect 404998 335696 405004 335708
rect 379440 335668 405004 335696
rect 379333 335659 379391 335665
rect 404998 335656 405004 335668
rect 405056 335656 405062 335708
rect 364794 335588 364800 335640
rect 364852 335628 364858 335640
rect 365530 335628 365536 335640
rect 364852 335600 365536 335628
rect 364852 335588 364858 335600
rect 365530 335588 365536 335600
rect 365588 335588 365594 335640
rect 368934 335588 368940 335640
rect 368992 335628 368998 335640
rect 370869 335631 370927 335637
rect 370869 335628 370881 335631
rect 368992 335600 370881 335628
rect 368992 335588 368998 335600
rect 370869 335597 370881 335600
rect 370915 335597 370927 335631
rect 398098 335628 398104 335640
rect 370869 335591 370927 335597
rect 370976 335600 398104 335628
rect 364306 335532 365300 335560
rect 193858 335452 193864 335504
rect 193916 335492 193922 335504
rect 266354 335492 266360 335504
rect 193916 335464 266360 335492
rect 193916 335452 193922 335464
rect 266354 335452 266360 335464
rect 266412 335452 266418 335504
rect 322290 335452 322296 335504
rect 322348 335492 322354 335504
rect 322842 335492 322848 335504
rect 322348 335464 322848 335492
rect 322348 335452 322354 335464
rect 322842 335452 322848 335464
rect 322900 335452 322906 335504
rect 327718 335492 327724 335504
rect 325666 335464 327724 335492
rect 191098 335384 191104 335436
rect 191156 335424 191162 335436
rect 265986 335424 265992 335436
rect 191156 335396 265992 335424
rect 191156 335384 191162 335396
rect 265986 335384 265992 335396
rect 266044 335384 266050 335436
rect 318978 335384 318984 335436
rect 319036 335424 319042 335436
rect 325666 335424 325694 335464
rect 327718 335452 327724 335464
rect 327776 335452 327782 335504
rect 363874 335452 363880 335504
rect 363932 335492 363938 335504
rect 364242 335492 364248 335504
rect 363932 335464 364248 335492
rect 363932 335452 363938 335464
rect 364242 335452 364248 335464
rect 364300 335452 364306 335504
rect 319036 335396 325694 335424
rect 319036 335384 319042 335396
rect 326522 335384 326528 335436
rect 326580 335424 326586 335436
rect 326890 335424 326896 335436
rect 326580 335396 326896 335424
rect 326580 335384 326586 335396
rect 326890 335384 326896 335396
rect 326948 335384 326954 335436
rect 336090 335384 336096 335436
rect 336148 335424 336154 335436
rect 336458 335424 336464 335436
rect 336148 335396 336464 335424
rect 336148 335384 336154 335396
rect 336458 335384 336464 335396
rect 336516 335384 336522 335436
rect 243538 335316 243544 335368
rect 243596 335356 243602 335368
rect 277394 335356 277400 335368
rect 243596 335328 277400 335356
rect 243596 335316 243602 335328
rect 277394 335316 277400 335328
rect 277452 335316 277458 335368
rect 315666 335316 315672 335368
rect 315724 335356 315730 335368
rect 317506 335356 317512 335368
rect 315724 335328 317512 335356
rect 315724 335316 315730 335328
rect 317506 335316 317512 335328
rect 317564 335316 317570 335368
rect 352190 335316 352196 335368
rect 352248 335356 352254 335368
rect 365272 335356 365300 335532
rect 365346 335520 365352 335572
rect 365404 335560 365410 335572
rect 370976 335560 371004 335600
rect 398098 335588 398104 335600
rect 398156 335588 398162 335640
rect 365404 335532 371004 335560
rect 371881 335563 371939 335569
rect 365404 335520 365410 335532
rect 371881 335529 371893 335563
rect 371927 335560 371939 335563
rect 377398 335560 377404 335572
rect 371927 335532 377404 335560
rect 371927 335529 371939 335532
rect 371881 335523 371939 335529
rect 377398 335520 377404 335532
rect 377456 335520 377462 335572
rect 377493 335563 377551 335569
rect 377493 335529 377505 335563
rect 377539 335560 377551 335563
rect 403618 335560 403624 335572
rect 377539 335532 403624 335560
rect 377539 335529 377551 335532
rect 377493 335523 377551 335529
rect 403618 335520 403624 335532
rect 403676 335520 403682 335572
rect 370869 335495 370927 335501
rect 370869 335461 370881 335495
rect 370915 335492 370927 335495
rect 399478 335492 399484 335504
rect 370915 335464 399484 335492
rect 370915 335461 370927 335464
rect 370869 335455 370927 335461
rect 399478 335452 399484 335464
rect 399536 335452 399542 335504
rect 371881 335427 371939 335433
rect 371881 335424 371893 335427
rect 369826 335396 371893 335424
rect 369826 335356 369854 335396
rect 371881 335393 371893 335396
rect 371927 335393 371939 335427
rect 371881 335387 371939 335393
rect 371970 335384 371976 335436
rect 372028 335424 372034 335436
rect 372522 335424 372528 335436
rect 372028 335396 372528 335424
rect 372028 335384 372034 335396
rect 372522 335384 372528 335396
rect 372580 335384 372586 335436
rect 372798 335384 372804 335436
rect 372856 335424 372862 335436
rect 373902 335424 373908 335436
rect 372856 335396 373908 335424
rect 372856 335384 372862 335396
rect 373902 335384 373908 335396
rect 373960 335384 373966 335436
rect 377030 335384 377036 335436
rect 377088 335424 377094 335436
rect 377088 335396 378272 335424
rect 377088 335384 377094 335396
rect 352248 335328 352880 335356
rect 365272 335328 369854 335356
rect 352248 335316 352254 335328
rect 352852 335220 352880 335328
rect 370406 335316 370412 335368
rect 370464 335356 370470 335368
rect 370866 335356 370872 335368
rect 370464 335328 370872 335356
rect 370464 335316 370470 335328
rect 370866 335316 370872 335328
rect 370924 335316 370930 335368
rect 370958 335316 370964 335368
rect 371016 335356 371022 335368
rect 371142 335356 371148 335368
rect 371016 335328 371148 335356
rect 371016 335316 371022 335328
rect 371142 335316 371148 335328
rect 371200 335316 371206 335368
rect 371602 335316 371608 335368
rect 371660 335356 371666 335368
rect 372154 335356 372160 335368
rect 371660 335328 372160 335356
rect 371660 335316 371666 335328
rect 372154 335316 372160 335328
rect 372212 335316 372218 335368
rect 373166 335316 373172 335368
rect 373224 335356 373230 335368
rect 373534 335356 373540 335368
rect 373224 335328 373540 335356
rect 373224 335316 373230 335328
rect 373534 335316 373540 335328
rect 373592 335316 373598 335368
rect 373626 335316 373632 335368
rect 373684 335356 373690 335368
rect 373810 335356 373816 335368
rect 373684 335328 373816 335356
rect 373684 335316 373690 335328
rect 373810 335316 373816 335328
rect 373868 335316 373874 335368
rect 374638 335316 374644 335368
rect 374696 335356 374702 335368
rect 375006 335356 375012 335368
rect 374696 335328 375012 335356
rect 374696 335316 374702 335328
rect 375006 335316 375012 335328
rect 375064 335316 375070 335368
rect 375098 335316 375104 335368
rect 375156 335356 375162 335368
rect 375282 335356 375288 335368
rect 375156 335328 375288 335356
rect 375156 335316 375162 335328
rect 375282 335316 375288 335328
rect 375340 335316 375346 335368
rect 375834 335316 375840 335368
rect 375892 335356 375898 335368
rect 376478 335356 376484 335368
rect 375892 335328 376484 335356
rect 375892 335316 375898 335328
rect 376478 335316 376484 335328
rect 376536 335316 376542 335368
rect 377306 335316 377312 335368
rect 377364 335356 377370 335368
rect 378042 335356 378048 335368
rect 377364 335328 378048 335356
rect 377364 335316 377370 335328
rect 378042 335316 378048 335328
rect 378100 335316 378106 335368
rect 378244 335356 378272 335396
rect 378502 335384 378508 335436
rect 378560 335424 378566 335436
rect 379238 335424 379244 335436
rect 378560 335396 379244 335424
rect 378560 335384 378566 335396
rect 379238 335384 379244 335396
rect 379296 335384 379302 335436
rect 379425 335427 379483 335433
rect 379425 335393 379437 335427
rect 379471 335424 379483 335427
rect 396718 335424 396724 335436
rect 379471 335396 396724 335424
rect 379471 335393 379483 335396
rect 379425 335387 379483 335393
rect 396718 335384 396724 335396
rect 396776 335384 396782 335436
rect 378244 335328 379008 335356
rect 378980 335288 379008 335328
rect 379054 335316 379060 335368
rect 379112 335356 379118 335368
rect 379330 335356 379336 335368
rect 379112 335328 379336 335356
rect 379112 335316 379118 335328
rect 379330 335316 379336 335328
rect 379388 335316 379394 335368
rect 380713 335359 380771 335365
rect 379440 335328 380296 335356
rect 379440 335288 379468 335328
rect 378980 335260 379468 335288
rect 380268 335288 380296 335328
rect 380713 335325 380725 335359
rect 380759 335354 380771 335359
rect 380759 335326 380793 335354
rect 380759 335325 380771 335326
rect 380713 335319 380771 335325
rect 380728 335288 380756 335319
rect 380268 335260 380756 335288
rect 353110 335220 353116 335232
rect 352852 335192 353116 335220
rect 353110 335180 353116 335192
rect 353168 335180 353174 335232
rect 261110 330760 261116 330812
rect 261168 330760 261174 330812
rect 272150 330760 272156 330812
rect 272208 330760 272214 330812
rect 261128 330608 261156 330760
rect 272168 330608 272196 330760
rect 332410 330624 332416 330676
rect 332468 330624 332474 330676
rect 261110 330556 261116 330608
rect 261168 330556 261174 330608
rect 272150 330556 272156 330608
rect 272208 330556 272214 330608
rect 309134 330556 309140 330608
rect 309192 330596 309198 330608
rect 310330 330596 310336 330608
rect 309192 330568 310336 330596
rect 309192 330556 309198 330568
rect 310330 330556 310336 330568
rect 310388 330556 310394 330608
rect 254118 330488 254124 330540
rect 254176 330528 254182 330540
rect 254946 330528 254952 330540
rect 254176 330500 254952 330528
rect 254176 330488 254182 330500
rect 254946 330488 254952 330500
rect 255004 330488 255010 330540
rect 256694 330488 256700 330540
rect 256752 330528 256758 330540
rect 257338 330528 257344 330540
rect 256752 330500 257344 330528
rect 256752 330488 256758 330500
rect 257338 330488 257344 330500
rect 257396 330488 257402 330540
rect 259730 330488 259736 330540
rect 259788 330528 259794 330540
rect 260650 330528 260656 330540
rect 259788 330500 260656 330528
rect 259788 330488 259794 330500
rect 260650 330488 260656 330500
rect 260708 330488 260714 330540
rect 261018 330488 261024 330540
rect 261076 330528 261082 330540
rect 261570 330528 261576 330540
rect 261076 330500 261576 330528
rect 261076 330488 261082 330500
rect 261570 330488 261576 330500
rect 261628 330488 261634 330540
rect 262490 330488 262496 330540
rect 262548 330528 262554 330540
rect 263318 330528 263324 330540
rect 262548 330500 263324 330528
rect 262548 330488 262554 330500
rect 263318 330488 263324 330500
rect 263376 330488 263382 330540
rect 265066 330488 265072 330540
rect 265124 330528 265130 330540
rect 265710 330528 265716 330540
rect 265124 330500 265716 330528
rect 265124 330488 265130 330500
rect 265710 330488 265716 330500
rect 265768 330488 265774 330540
rect 266446 330488 266452 330540
rect 266504 330528 266510 330540
rect 266906 330528 266912 330540
rect 266504 330500 266912 330528
rect 266504 330488 266510 330500
rect 266906 330488 266912 330500
rect 266964 330488 266970 330540
rect 267918 330488 267924 330540
rect 267976 330528 267982 330540
rect 268746 330528 268752 330540
rect 267976 330500 268752 330528
rect 267976 330488 267982 330500
rect 268746 330488 268752 330500
rect 268804 330488 268810 330540
rect 269114 330488 269120 330540
rect 269172 330528 269178 330540
rect 269574 330528 269580 330540
rect 269172 330500 269580 330528
rect 269172 330488 269178 330500
rect 269574 330488 269580 330500
rect 269632 330488 269638 330540
rect 270770 330488 270776 330540
rect 270828 330528 270834 330540
rect 271690 330528 271696 330540
rect 270828 330500 271696 330528
rect 270828 330488 270834 330500
rect 271690 330488 271696 330500
rect 271748 330488 271754 330540
rect 272058 330488 272064 330540
rect 272116 330528 272122 330540
rect 272610 330528 272616 330540
rect 272116 330500 272616 330528
rect 272116 330488 272122 330500
rect 272610 330488 272616 330500
rect 272668 330488 272674 330540
rect 302418 330488 302424 330540
rect 302476 330528 302482 330540
rect 303430 330528 303436 330540
rect 302476 330500 303436 330528
rect 302476 330488 302482 330500
rect 303430 330488 303436 330500
rect 303488 330488 303494 330540
rect 305178 330488 305184 330540
rect 305236 330528 305242 330540
rect 305822 330528 305828 330540
rect 305236 330500 305828 330528
rect 305236 330488 305242 330500
rect 305822 330488 305828 330500
rect 305880 330488 305886 330540
rect 307846 330488 307852 330540
rect 307904 330528 307910 330540
rect 308490 330528 308496 330540
rect 307904 330500 308496 330528
rect 307904 330488 307910 330500
rect 308490 330488 308496 330500
rect 308548 330488 308554 330540
rect 309226 330488 309232 330540
rect 309284 330528 309290 330540
rect 309686 330528 309692 330540
rect 309284 330500 309692 330528
rect 309284 330488 309290 330500
rect 309686 330488 309692 330500
rect 309744 330488 309750 330540
rect 313274 330488 313280 330540
rect 313332 330528 313338 330540
rect 314194 330528 314200 330540
rect 313332 330500 314200 330528
rect 313332 330488 313338 330500
rect 314194 330488 314200 330500
rect 314252 330488 314258 330540
rect 266538 330420 266544 330472
rect 266596 330460 266602 330472
rect 267182 330460 267188 330472
rect 266596 330432 267188 330460
rect 266596 330420 266602 330432
rect 267182 330420 267188 330432
rect 267240 330420 267246 330472
rect 267734 330420 267740 330472
rect 267792 330460 267798 330472
rect 268378 330460 268384 330472
rect 267792 330432 268384 330460
rect 267792 330420 267798 330432
rect 268378 330420 268384 330432
rect 268436 330420 268442 330472
rect 269206 330420 269212 330472
rect 269264 330460 269270 330472
rect 269942 330460 269948 330472
rect 269264 330432 269948 330460
rect 269264 330420 269270 330432
rect 269942 330420 269948 330432
rect 270000 330420 270006 330472
rect 270586 330420 270592 330472
rect 270644 330460 270650 330472
rect 271414 330460 271420 330472
rect 270644 330432 271420 330460
rect 270644 330420 270650 330432
rect 271414 330420 271420 330432
rect 271472 330420 271478 330472
rect 271874 330420 271880 330472
rect 271932 330460 271938 330472
rect 272886 330460 272892 330472
rect 271932 330432 272892 330460
rect 271932 330420 271938 330432
rect 272886 330420 272892 330432
rect 272944 330420 272950 330472
rect 307938 330420 307944 330472
rect 307996 330460 308002 330472
rect 308766 330460 308772 330472
rect 307996 330432 308772 330460
rect 307996 330420 308002 330432
rect 308766 330420 308772 330432
rect 308824 330420 308830 330472
rect 309318 330420 309324 330472
rect 309376 330460 309382 330472
rect 309962 330460 309968 330472
rect 309376 330432 309968 330460
rect 309376 330420 309382 330432
rect 309962 330420 309968 330432
rect 310020 330420 310026 330472
rect 320450 330420 320456 330472
rect 320508 330460 320514 330472
rect 321370 330460 321376 330472
rect 320508 330432 321376 330460
rect 320508 330420 320514 330432
rect 321370 330420 321376 330432
rect 321428 330420 321434 330472
rect 323762 330420 323768 330472
rect 323820 330460 323826 330472
rect 324038 330460 324044 330472
rect 323820 330432 324044 330460
rect 323820 330420 323826 330432
rect 324038 330420 324044 330432
rect 324096 330420 324102 330472
rect 326154 330420 326160 330472
rect 326212 330460 326218 330472
rect 326706 330460 326712 330472
rect 326212 330432 326712 330460
rect 326212 330420 326218 330432
rect 326706 330420 326712 330432
rect 326764 330420 326770 330472
rect 332226 330420 332232 330472
rect 332284 330460 332290 330472
rect 332428 330460 332456 330624
rect 370130 330488 370136 330540
rect 370188 330528 370194 330540
rect 371050 330528 371056 330540
rect 370188 330500 371056 330528
rect 370188 330488 370194 330500
rect 371050 330488 371056 330500
rect 371108 330488 371114 330540
rect 374362 330488 374368 330540
rect 374420 330528 374426 330540
rect 375190 330528 375196 330540
rect 374420 330500 375196 330528
rect 374420 330488 374426 330500
rect 375190 330488 375196 330500
rect 375248 330488 375254 330540
rect 376386 330488 376392 330540
rect 376444 330528 376450 330540
rect 376662 330528 376668 330540
rect 376444 330500 376668 330528
rect 376444 330488 376450 330500
rect 376662 330488 376668 330500
rect 376720 330488 376726 330540
rect 332284 330432 332456 330460
rect 332284 330420 332290 330432
rect 357158 330420 357164 330472
rect 357216 330460 357222 330472
rect 357434 330460 357440 330472
rect 357216 330432 357440 330460
rect 357216 330420 357222 330432
rect 357434 330420 357440 330432
rect 357492 330420 357498 330472
rect 302326 328924 302332 328976
rect 302384 328964 302390 328976
rect 303154 328964 303160 328976
rect 302384 328936 303160 328964
rect 302384 328924 302390 328936
rect 303154 328924 303160 328936
rect 303212 328924 303218 328976
rect 255406 327632 255412 327684
rect 255464 327672 255470 327684
rect 256142 327672 256148 327684
rect 255464 327644 256148 327672
rect 255464 327632 255470 327644
rect 256142 327632 256148 327644
rect 256200 327632 256206 327684
rect 288710 326816 288716 326868
rect 288768 326816 288774 326868
rect 256878 326748 256884 326800
rect 256936 326788 256942 326800
rect 257614 326788 257620 326800
rect 256936 326760 257620 326788
rect 256936 326748 256942 326760
rect 257614 326748 257620 326760
rect 257672 326748 257678 326800
rect 278774 326680 278780 326732
rect 278832 326720 278838 326732
rect 279050 326720 279056 326732
rect 278832 326692 279056 326720
rect 278832 326680 278838 326692
rect 279050 326680 279056 326692
rect 279108 326680 279114 326732
rect 284478 326680 284484 326732
rect 284536 326720 284542 326732
rect 284754 326720 284760 326732
rect 284536 326692 284760 326720
rect 284536 326680 284542 326692
rect 284754 326680 284760 326692
rect 284812 326680 284818 326732
rect 288728 326664 288756 326816
rect 293862 326680 293868 326732
rect 293920 326720 293926 326732
rect 294414 326720 294420 326732
rect 293920 326692 294420 326720
rect 293920 326680 293926 326692
rect 294414 326680 294420 326692
rect 294472 326680 294478 326732
rect 288710 326612 288716 326664
rect 288768 326612 288774 326664
rect 262398 326544 262404 326596
rect 262456 326584 262462 326596
rect 263042 326584 263048 326596
rect 262456 326556 263048 326584
rect 262456 326544 262462 326556
rect 263042 326544 263048 326556
rect 263100 326544 263106 326596
rect 287054 326476 287060 326528
rect 287112 326516 287118 326528
rect 287330 326516 287336 326528
rect 287112 326488 287336 326516
rect 287112 326476 287118 326488
rect 287330 326476 287336 326488
rect 287388 326476 287394 326528
rect 294046 326476 294052 326528
rect 294104 326516 294110 326528
rect 294322 326516 294328 326528
rect 294104 326488 294328 326516
rect 294104 326476 294110 326488
rect 294322 326476 294328 326488
rect 294380 326476 294386 326528
rect 295518 326516 295524 326528
rect 295479 326488 295524 326516
rect 295518 326476 295524 326488
rect 295576 326476 295582 326528
rect 244550 326408 244556 326460
rect 244608 326448 244614 326460
rect 245102 326448 245108 326460
rect 244608 326420 245108 326448
rect 244608 326408 244614 326420
rect 245102 326408 245108 326420
rect 245160 326408 245166 326460
rect 245930 326408 245936 326460
rect 245988 326448 245994 326460
rect 246574 326448 246580 326460
rect 245988 326420 246580 326448
rect 245988 326408 245994 326420
rect 246574 326408 246580 326420
rect 246632 326408 246638 326460
rect 247310 326408 247316 326460
rect 247368 326448 247374 326460
rect 248046 326448 248052 326460
rect 247368 326420 248052 326448
rect 247368 326408 247374 326420
rect 248046 326408 248052 326420
rect 248104 326408 248110 326460
rect 252738 326408 252744 326460
rect 252796 326448 252802 326460
rect 253474 326448 253480 326460
rect 252796 326420 253480 326448
rect 252796 326408 252802 326420
rect 253474 326408 253480 326420
rect 253532 326408 253538 326460
rect 276198 326408 276204 326460
rect 276256 326448 276262 326460
rect 277118 326448 277124 326460
rect 276256 326420 277124 326448
rect 276256 326408 276262 326420
rect 277118 326408 277124 326420
rect 277176 326408 277182 326460
rect 280246 326408 280252 326460
rect 280304 326448 280310 326460
rect 280982 326448 280988 326460
rect 280304 326420 280988 326448
rect 280304 326408 280310 326420
rect 280982 326408 280988 326420
rect 281040 326408 281046 326460
rect 281718 326408 281724 326460
rect 281776 326448 281782 326460
rect 282454 326448 282460 326460
rect 281776 326420 282460 326448
rect 281776 326408 281782 326420
rect 282454 326408 282460 326420
rect 282512 326408 282518 326460
rect 283098 326408 283104 326460
rect 283156 326448 283162 326460
rect 283926 326448 283932 326460
rect 283156 326420 283932 326448
rect 283156 326408 283162 326420
rect 283926 326408 283932 326420
rect 283984 326408 283990 326460
rect 284386 326408 284392 326460
rect 284444 326448 284450 326460
rect 285490 326448 285496 326460
rect 284444 326420 285496 326448
rect 284444 326408 284450 326420
rect 285490 326408 285496 326420
rect 285548 326408 285554 326460
rect 288434 326408 288440 326460
rect 288492 326448 288498 326460
rect 289078 326448 289084 326460
rect 288492 326420 289084 326448
rect 288492 326408 288498 326420
rect 289078 326408 289084 326420
rect 289136 326408 289142 326460
rect 291194 326408 291200 326460
rect 291252 326448 291258 326460
rect 291746 326448 291752 326460
rect 291252 326420 291752 326448
rect 291252 326408 291258 326420
rect 291746 326408 291752 326420
rect 291804 326408 291810 326460
rect 296898 326408 296904 326460
rect 296956 326448 296962 326460
rect 297726 326448 297732 326460
rect 296956 326420 297732 326448
rect 296956 326408 296962 326420
rect 297726 326408 297732 326420
rect 297784 326408 297790 326460
rect 234706 326340 234712 326392
rect 234764 326380 234770 326392
rect 235534 326380 235540 326392
rect 234764 326352 235540 326380
rect 234764 326340 234770 326352
rect 235534 326340 235540 326352
rect 235592 326340 235598 326392
rect 236086 326340 236092 326392
rect 236144 326380 236150 326392
rect 236730 326380 236736 326392
rect 236144 326352 236736 326380
rect 236144 326340 236150 326352
rect 236730 326340 236736 326352
rect 236788 326340 236794 326392
rect 237374 326340 237380 326392
rect 237432 326380 237438 326392
rect 238478 326380 238484 326392
rect 237432 326352 238484 326380
rect 237432 326340 237438 326352
rect 238478 326340 238484 326352
rect 238536 326340 238542 326392
rect 238846 326340 238852 326392
rect 238904 326380 238910 326392
rect 239674 326380 239680 326392
rect 238904 326352 239680 326380
rect 238904 326340 238910 326352
rect 239674 326340 239680 326352
rect 239732 326340 239738 326392
rect 240318 326340 240324 326392
rect 240376 326380 240382 326392
rect 240870 326380 240876 326392
rect 240376 326352 240876 326380
rect 240376 326340 240382 326352
rect 240870 326340 240876 326352
rect 240928 326340 240934 326392
rect 241606 326340 241612 326392
rect 241664 326380 241670 326392
rect 242066 326380 242072 326392
rect 241664 326352 242072 326380
rect 241664 326340 241670 326352
rect 242066 326340 242072 326352
rect 242124 326340 242130 326392
rect 244366 326340 244372 326392
rect 244424 326380 244430 326392
rect 244826 326380 244832 326392
rect 244424 326352 244832 326380
rect 244424 326340 244430 326352
rect 244826 326340 244832 326352
rect 244884 326340 244890 326392
rect 245746 326340 245752 326392
rect 245804 326380 245810 326392
rect 246298 326380 246304 326392
rect 245804 326352 246304 326380
rect 245804 326340 245810 326352
rect 246298 326340 246304 326352
rect 246356 326340 246362 326392
rect 247218 326340 247224 326392
rect 247276 326380 247282 326392
rect 247770 326380 247776 326392
rect 247276 326352 247776 326380
rect 247276 326340 247282 326352
rect 247770 326340 247776 326352
rect 247828 326340 247834 326392
rect 248506 326340 248512 326392
rect 248564 326380 248570 326392
rect 249610 326380 249616 326392
rect 248564 326352 249616 326380
rect 248564 326340 248570 326352
rect 249610 326340 249616 326352
rect 249668 326340 249674 326392
rect 249886 326340 249892 326392
rect 249944 326380 249950 326392
rect 250806 326380 250812 326392
rect 249944 326352 250812 326380
rect 249944 326340 249950 326352
rect 250806 326340 250812 326352
rect 250864 326340 250870 326392
rect 251266 326340 251272 326392
rect 251324 326380 251330 326392
rect 252278 326380 252284 326392
rect 251324 326352 252284 326380
rect 251324 326340 251330 326352
rect 252278 326340 252284 326352
rect 252336 326340 252342 326392
rect 252646 326340 252652 326392
rect 252704 326380 252710 326392
rect 253198 326380 253204 326392
rect 252704 326352 253204 326380
rect 252704 326340 252710 326352
rect 253198 326340 253204 326352
rect 253256 326340 253262 326392
rect 273438 326340 273444 326392
rect 273496 326380 273502 326392
rect 274082 326380 274088 326392
rect 273496 326352 274088 326380
rect 273496 326340 273502 326352
rect 274082 326340 274088 326352
rect 274140 326340 274146 326392
rect 276106 326340 276112 326392
rect 276164 326380 276170 326392
rect 276750 326380 276756 326392
rect 276164 326352 276756 326380
rect 276164 326340 276170 326352
rect 276750 326340 276756 326352
rect 276808 326340 276814 326392
rect 278866 326340 278872 326392
rect 278924 326380 278930 326392
rect 279510 326380 279516 326392
rect 278924 326352 279516 326380
rect 278924 326340 278930 326352
rect 279510 326340 279516 326352
rect 279568 326340 279574 326392
rect 280430 326340 280436 326392
rect 280488 326380 280494 326392
rect 281258 326380 281264 326392
rect 280488 326352 281264 326380
rect 280488 326340 280494 326352
rect 281258 326340 281264 326352
rect 281316 326340 281322 326392
rect 281626 326340 281632 326392
rect 281684 326380 281690 326392
rect 282178 326380 282184 326392
rect 281684 326352 282184 326380
rect 281684 326340 281690 326352
rect 282178 326340 282184 326352
rect 282236 326340 282242 326392
rect 283006 326340 283012 326392
rect 283064 326380 283070 326392
rect 283650 326380 283656 326392
rect 283064 326352 283656 326380
rect 283064 326340 283070 326352
rect 283650 326340 283656 326352
rect 283708 326340 283714 326392
rect 284570 326340 284576 326392
rect 284628 326380 284634 326392
rect 285214 326380 285220 326392
rect 284628 326352 285220 326380
rect 284628 326340 284634 326352
rect 285214 326340 285220 326352
rect 285272 326340 285278 326392
rect 287330 326340 287336 326392
rect 287388 326380 287394 326392
rect 287882 326380 287888 326392
rect 287388 326352 287888 326380
rect 287388 326340 287394 326352
rect 287882 326340 287888 326352
rect 287940 326340 287946 326392
rect 288618 326340 288624 326392
rect 288676 326380 288682 326392
rect 289354 326380 289360 326392
rect 288676 326352 289360 326380
rect 288676 326340 288682 326352
rect 289354 326340 289360 326352
rect 289412 326340 289418 326392
rect 289906 326340 289912 326392
rect 289964 326380 289970 326392
rect 290550 326380 290556 326392
rect 289964 326352 290556 326380
rect 289964 326340 289970 326352
rect 290550 326340 290556 326352
rect 290608 326340 290614 326392
rect 291470 326340 291476 326392
rect 291528 326380 291534 326392
rect 292390 326380 292396 326392
rect 291528 326352 292396 326380
rect 291528 326340 291534 326352
rect 292390 326340 292396 326352
rect 292448 326340 292454 326392
rect 296806 326340 296812 326392
rect 296864 326380 296870 326392
rect 297450 326380 297456 326392
rect 296864 326352 297456 326380
rect 296864 326340 296870 326352
rect 297450 326340 297456 326352
rect 297508 326340 297514 326392
rect 298278 326340 298284 326392
rect 298336 326380 298342 326392
rect 299198 326380 299204 326392
rect 298336 326352 299204 326380
rect 298336 326340 298342 326352
rect 299198 326340 299204 326352
rect 299256 326340 299262 326392
rect 299566 326340 299572 326392
rect 299624 326380 299630 326392
rect 300118 326380 300124 326392
rect 299624 326352 300124 326380
rect 299624 326340 299630 326352
rect 300118 326340 300124 326352
rect 300176 326340 300182 326392
rect 247034 326272 247040 326324
rect 247092 326312 247098 326324
rect 247494 326312 247500 326324
rect 247092 326284 247500 326312
rect 247092 326272 247098 326284
rect 247494 326272 247500 326284
rect 247552 326272 247558 326324
rect 291286 326272 291292 326324
rect 291344 326312 291350 326324
rect 292022 326312 292028 326324
rect 291344 326284 292028 326312
rect 291344 326272 291350 326284
rect 292022 326272 292028 326284
rect 292080 326272 292086 326324
rect 292574 324232 292580 324284
rect 292632 324272 292638 324284
rect 293586 324272 293592 324284
rect 292632 324244 293592 324272
rect 292632 324232 292638 324244
rect 293586 324232 293592 324244
rect 293644 324232 293650 324284
rect 242986 323552 242992 323604
rect 243044 323592 243050 323604
rect 243170 323592 243176 323604
rect 243044 323564 243176 323592
rect 243044 323552 243050 323564
rect 243170 323552 243176 323564
rect 243228 323552 243234 323604
rect 285674 323552 285680 323604
rect 285732 323592 285738 323604
rect 286410 323592 286416 323604
rect 285732 323564 286416 323592
rect 285732 323552 285738 323564
rect 286410 323552 286416 323564
rect 286468 323552 286474 323604
rect 288526 323552 288532 323604
rect 288584 323592 288590 323604
rect 288802 323592 288808 323604
rect 288584 323564 288808 323592
rect 288584 323552 288590 323564
rect 288802 323552 288808 323564
rect 288860 323552 288866 323604
rect 295518 323592 295524 323604
rect 295479 323564 295524 323592
rect 295518 323552 295524 323564
rect 295576 323552 295582 323604
rect 273254 323280 273260 323332
rect 273312 323320 273318 323332
rect 273806 323320 273812 323332
rect 273312 323292 273812 323320
rect 273312 323280 273318 323292
rect 273806 323280 273812 323292
rect 273864 323280 273870 323332
rect 236178 323144 236184 323196
rect 236236 323184 236242 323196
rect 237006 323184 237012 323196
rect 236236 323156 237012 323184
rect 236236 323144 236242 323156
rect 237006 323144 237012 323156
rect 237064 323144 237070 323196
rect 240226 321852 240232 321904
rect 240284 321892 240290 321904
rect 240594 321892 240600 321904
rect 240284 321864 240600 321892
rect 240284 321852 240290 321864
rect 240594 321852 240600 321864
rect 240652 321852 240658 321904
rect 287146 321784 287152 321836
rect 287204 321824 287210 321836
rect 288158 321824 288164 321836
rect 287204 321796 288164 321824
rect 287204 321784 287210 321796
rect 288158 321784 288164 321796
rect 288216 321784 288222 321836
rect 251450 320696 251456 320748
rect 251508 320736 251514 320748
rect 251634 320736 251640 320748
rect 251508 320708 251640 320736
rect 251508 320696 251514 320708
rect 251634 320696 251640 320708
rect 251692 320696 251698 320748
rect 2774 319812 2780 319864
rect 2832 319852 2838 319864
rect 5166 319852 5172 319864
rect 2832 319824 5172 319852
rect 2832 319812 2838 319824
rect 5166 319812 5172 319824
rect 5224 319812 5230 319864
rect 238938 319540 238944 319592
rect 238996 319580 239002 319592
rect 239122 319580 239128 319592
rect 238996 319552 239128 319580
rect 238996 319540 239002 319552
rect 239122 319540 239128 319552
rect 239180 319540 239186 319592
rect 383562 299412 383568 299464
rect 383620 299452 383626 299464
rect 580166 299452 580172 299464
rect 383620 299424 580172 299452
rect 383620 299412 383626 299424
rect 580166 299412 580172 299424
rect 580224 299412 580230 299464
rect 3142 293768 3148 293820
rect 3200 293808 3206 293820
rect 6546 293808 6552 293820
rect 3200 293780 6552 293808
rect 3200 293768 3206 293780
rect 6546 293768 6552 293780
rect 6604 293768 6610 293820
rect 385770 273164 385776 273216
rect 385828 273204 385834 273216
rect 580166 273204 580172 273216
rect 385828 273176 580172 273204
rect 385828 273164 385834 273176
rect 580166 273164 580172 273176
rect 580224 273164 580230 273216
rect 2774 267248 2780 267300
rect 2832 267288 2838 267300
rect 5074 267288 5080 267300
rect 2832 267260 5080 267288
rect 2832 267248 2838 267260
rect 5074 267248 5080 267260
rect 5132 267248 5138 267300
rect 383470 245556 383476 245608
rect 383528 245596 383534 245608
rect 580166 245596 580172 245608
rect 383528 245568 580172 245596
rect 383528 245556 383534 245568
rect 580166 245556 580172 245568
rect 580224 245556 580230 245608
rect 3234 241068 3240 241120
rect 3292 241108 3298 241120
rect 6454 241108 6460 241120
rect 3292 241080 6460 241108
rect 3292 241068 3298 241080
rect 6454 241068 6460 241080
rect 6512 241068 6518 241120
rect 384850 233180 384856 233232
rect 384908 233220 384914 233232
rect 579982 233220 579988 233232
rect 384908 233192 579988 233220
rect 384908 233180 384914 233192
rect 579982 233180 579988 233192
rect 580040 233180 580046 233232
rect 383378 206932 383384 206984
rect 383436 206972 383442 206984
rect 580166 206972 580172 206984
rect 383436 206944 580172 206972
rect 383436 206932 383442 206944
rect 580166 206932 580172 206944
rect 580224 206932 580230 206984
rect 384758 193128 384764 193180
rect 384816 193168 384822 193180
rect 580166 193168 580172 193180
rect 384816 193140 580172 193168
rect 384816 193128 384822 193140
rect 580166 193128 580172 193140
rect 580224 193128 580230 193180
rect 3234 188844 3240 188896
rect 3292 188884 3298 188896
rect 6362 188884 6368 188896
rect 3292 188856 6368 188884
rect 3292 188844 3298 188856
rect 6362 188844 6368 188856
rect 6420 188844 6426 188896
rect 383286 166948 383292 167000
rect 383344 166988 383350 167000
rect 580166 166988 580172 167000
rect 383344 166960 580172 166988
rect 383344 166948 383350 166960
rect 580166 166948 580172 166960
rect 580224 166948 580230 167000
rect 384666 153144 384672 153196
rect 384724 153184 384730 153196
rect 579614 153184 579620 153196
rect 384724 153156 579620 153184
rect 384724 153144 384730 153156
rect 579614 153144 579620 153156
rect 579672 153144 579678 153196
rect 3234 137844 3240 137896
rect 3292 137884 3298 137896
rect 6270 137884 6276 137896
rect 3292 137856 6276 137884
rect 3292 137844 3298 137856
rect 6270 137844 6276 137856
rect 6328 137844 6334 137896
rect 383102 126896 383108 126948
rect 383160 126936 383166 126948
rect 580166 126936 580172 126948
rect 383160 126908 580172 126936
rect 383160 126896 383166 126908
rect 580166 126896 580172 126908
rect 580224 126896 580230 126948
rect 384574 113092 384580 113144
rect 384632 113132 384638 113144
rect 580166 113132 580172 113144
rect 384632 113104 580172 113132
rect 384632 113092 384638 113104
rect 580166 113092 580172 113104
rect 580224 113092 580230 113144
rect 2774 110712 2780 110764
rect 2832 110752 2838 110764
rect 4982 110752 4988 110764
rect 2832 110724 4988 110752
rect 2832 110712 2838 110724
rect 4982 110712 4988 110724
rect 5040 110712 5046 110764
rect 3326 97860 3332 97912
rect 3384 97900 3390 97912
rect 8018 97900 8024 97912
rect 3384 97872 8024 97900
rect 3384 97860 3390 97872
rect 8018 97860 8024 97872
rect 8076 97860 8082 97912
rect 383010 86912 383016 86964
rect 383068 86952 383074 86964
rect 580166 86952 580172 86964
rect 383068 86924 580172 86952
rect 383068 86912 383074 86924
rect 580166 86912 580172 86924
rect 580224 86912 580230 86964
rect 2774 85008 2780 85060
rect 2832 85048 2838 85060
rect 6178 85048 6184 85060
rect 2832 85020 6184 85048
rect 2832 85008 2838 85020
rect 6178 85008 6184 85020
rect 6236 85008 6242 85060
rect 384390 73108 384396 73160
rect 384448 73148 384454 73160
rect 580166 73148 580172 73160
rect 384448 73120 580172 73148
rect 384448 73108 384454 73120
rect 580166 73108 580172 73120
rect 580224 73108 580230 73160
rect 2774 71612 2780 71664
rect 2832 71652 2838 71664
rect 4890 71652 4896 71664
rect 2832 71624 4896 71652
rect 2832 71612 2838 71624
rect 4890 71612 4896 71624
rect 4948 71612 4954 71664
rect 385678 60664 385684 60716
rect 385736 60704 385742 60716
rect 580166 60704 580172 60716
rect 385736 60676 580172 60704
rect 385736 60664 385742 60676
rect 580166 60664 580172 60676
rect 580224 60664 580230 60716
rect 3050 59304 3056 59356
rect 3108 59344 3114 59356
rect 7834 59344 7840 59356
rect 3108 59316 7840 59344
rect 3108 59304 3114 59316
rect 7834 59304 7840 59316
rect 7892 59304 7898 59356
rect 382918 46860 382924 46912
rect 382976 46900 382982 46912
rect 580166 46900 580172 46912
rect 382976 46872 580172 46900
rect 382976 46860 382982 46872
rect 580166 46860 580172 46872
rect 580224 46860 580230 46912
rect 3418 45500 3424 45552
rect 3476 45540 3482 45552
rect 7742 45540 7748 45552
rect 3476 45512 7748 45540
rect 3476 45500 3482 45512
rect 7742 45500 7748 45512
rect 7800 45500 7806 45552
rect 384482 33056 384488 33108
rect 384540 33096 384546 33108
rect 580166 33096 580172 33108
rect 384540 33068 580172 33096
rect 384540 33056 384546 33068
rect 580166 33056 580172 33068
rect 580224 33056 580230 33108
rect 2774 32988 2780 33040
rect 2832 33028 2838 33040
rect 4798 33028 4804 33040
rect 2832 33000 4804 33028
rect 2832 32988 2838 33000
rect 4798 32988 4804 33000
rect 4856 32988 4862 33040
rect 384298 20612 384304 20664
rect 384356 20652 384362 20664
rect 579982 20652 579988 20664
rect 384356 20624 579988 20652
rect 384356 20612 384362 20624
rect 579982 20612 579988 20624
rect 580040 20612 580046 20664
rect 3050 20136 3056 20188
rect 3108 20176 3114 20188
rect 7650 20176 7656 20188
rect 3108 20148 7656 20176
rect 3108 20136 3114 20148
rect 7650 20136 7656 20148
rect 7708 20136 7714 20188
rect 119890 13472 119896 13524
rect 119948 13512 119954 13524
rect 265158 13512 265164 13524
rect 119948 13484 265164 13512
rect 119948 13472 119954 13484
rect 265158 13472 265164 13484
rect 265216 13472 265222 13524
rect 117222 13404 117228 13456
rect 117280 13444 117286 13456
rect 263778 13444 263784 13456
rect 117280 13416 263784 13444
rect 117280 13404 117286 13416
rect 263778 13404 263784 13416
rect 263836 13404 263842 13456
rect 112806 13336 112812 13388
rect 112864 13376 112870 13388
rect 262490 13376 262496 13388
rect 112864 13348 262496 13376
rect 112864 13336 112870 13348
rect 262490 13336 262496 13348
rect 262548 13336 262554 13388
rect 110322 13268 110328 13320
rect 110380 13308 110386 13320
rect 262582 13308 262588 13320
rect 110380 13280 262588 13308
rect 110380 13268 110386 13280
rect 262582 13268 262588 13280
rect 262640 13268 262646 13320
rect 106182 13200 106188 13252
rect 106240 13240 106246 13252
rect 261018 13240 261024 13252
rect 106240 13212 261024 13240
rect 106240 13200 106246 13212
rect 261018 13200 261024 13212
rect 261076 13200 261082 13252
rect 103422 13132 103428 13184
rect 103480 13172 103486 13184
rect 259730 13172 259736 13184
rect 103480 13144 259736 13172
rect 103480 13132 103486 13144
rect 259730 13132 259736 13144
rect 259788 13132 259794 13184
rect 99282 13064 99288 13116
rect 99340 13104 99346 13116
rect 259638 13104 259644 13116
rect 99340 13076 259644 13104
rect 99340 13064 99346 13076
rect 259638 13064 259644 13076
rect 259696 13064 259702 13116
rect 248414 12520 248420 12572
rect 248472 12560 248478 12572
rect 248690 12560 248696 12572
rect 248472 12532 248696 12560
rect 248472 12520 248478 12532
rect 248690 12520 248696 12532
rect 248748 12520 248754 12572
rect 161290 12384 161296 12436
rect 161348 12424 161354 12436
rect 274910 12424 274916 12436
rect 161348 12396 274916 12424
rect 161348 12384 161354 12396
rect 274910 12384 274916 12396
rect 274968 12384 274974 12436
rect 160094 12316 160100 12368
rect 160152 12356 160158 12368
rect 274818 12356 274824 12368
rect 160152 12328 274824 12356
rect 160152 12316 160158 12328
rect 274818 12316 274824 12328
rect 274876 12316 274882 12368
rect 147582 12248 147588 12300
rect 147640 12288 147646 12300
rect 272150 12288 272156 12300
rect 147640 12260 272156 12288
rect 147640 12248 147646 12260
rect 272150 12248 272156 12260
rect 272208 12248 272214 12300
rect 144822 12180 144828 12232
rect 144880 12220 144886 12232
rect 270862 12220 270868 12232
rect 144880 12192 270868 12220
rect 144880 12180 144886 12192
rect 270862 12180 270868 12192
rect 270920 12180 270926 12232
rect 362494 12180 362500 12232
rect 362552 12220 362558 12232
rect 503714 12220 503720 12232
rect 362552 12192 503720 12220
rect 362552 12180 362558 12192
rect 503714 12180 503720 12192
rect 503772 12180 503778 12232
rect 140038 12112 140044 12164
rect 140096 12152 140102 12164
rect 269482 12152 269488 12164
rect 140096 12124 269488 12152
rect 140096 12112 140102 12124
rect 269482 12112 269488 12124
rect 269540 12112 269546 12164
rect 363966 12112 363972 12164
rect 364024 12152 364030 12164
rect 507210 12152 507216 12164
rect 364024 12124 507216 12152
rect 364024 12112 364030 12124
rect 507210 12112 507216 12124
rect 507268 12112 507274 12164
rect 136450 12044 136456 12096
rect 136508 12084 136514 12096
rect 269390 12084 269396 12096
rect 136508 12056 269396 12084
rect 136508 12044 136514 12056
rect 269390 12044 269396 12056
rect 269448 12044 269454 12096
rect 366726 12044 366732 12096
rect 366784 12084 366790 12096
rect 517882 12084 517888 12096
rect 366784 12056 517888 12084
rect 366784 12044 366790 12056
rect 517882 12044 517888 12056
rect 517940 12044 517946 12096
rect 125870 11976 125876 12028
rect 125928 12016 125934 12028
rect 266630 12016 266636 12028
rect 125928 11988 266636 12016
rect 125928 11976 125934 11988
rect 266630 11976 266636 11988
rect 266688 11976 266694 12028
rect 368106 11976 368112 12028
rect 368164 12016 368170 12028
rect 525426 12016 525432 12028
rect 368164 11988 525432 12016
rect 368164 11976 368170 11988
rect 525426 11976 525432 11988
rect 525484 11976 525490 12028
rect 95142 11908 95148 11960
rect 95200 11948 95206 11960
rect 258350 11948 258356 11960
rect 95200 11920 258356 11948
rect 95200 11908 95206 11920
rect 258350 11908 258356 11920
rect 258408 11908 258414 11960
rect 372338 11908 372344 11960
rect 372396 11948 372402 11960
rect 539594 11948 539600 11960
rect 372396 11920 539600 11948
rect 372396 11908 372402 11920
rect 539594 11908 539600 11920
rect 539652 11908 539658 11960
rect 92382 11840 92388 11892
rect 92440 11880 92446 11892
rect 258258 11880 258264 11892
rect 92440 11852 258264 11880
rect 92440 11840 92446 11852
rect 258258 11840 258264 11852
rect 258316 11840 258322 11892
rect 373534 11840 373540 11892
rect 373592 11880 373598 11892
rect 546678 11880 546684 11892
rect 373592 11852 546684 11880
rect 373592 11840 373598 11852
rect 546678 11840 546684 11852
rect 546736 11840 546742 11892
rect 87966 11772 87972 11824
rect 88024 11812 88030 11824
rect 256970 11812 256976 11824
rect 88024 11784 256976 11812
rect 88024 11772 88030 11784
rect 256970 11772 256976 11784
rect 257028 11772 257034 11824
rect 380526 11772 380532 11824
rect 380584 11812 380590 11824
rect 575106 11812 575112 11824
rect 380584 11784 575112 11812
rect 380584 11772 380590 11784
rect 575106 11772 575112 11784
rect 575164 11772 575170 11824
rect 85482 11704 85488 11756
rect 85540 11744 85546 11756
rect 255406 11744 255412 11756
rect 85540 11716 255412 11744
rect 85540 11704 85546 11716
rect 255406 11704 255412 11716
rect 255464 11704 255470 11756
rect 381998 11704 382004 11756
rect 382056 11744 382062 11756
rect 580994 11744 581000 11756
rect 382056 11716 581000 11744
rect 382056 11704 382062 11716
rect 580994 11704 581000 11716
rect 581052 11704 581058 11756
rect 164878 11636 164884 11688
rect 164936 11676 164942 11688
rect 276382 11676 276388 11688
rect 164936 11648 276388 11676
rect 164936 11636 164942 11648
rect 276382 11636 276388 11648
rect 276440 11636 276446 11688
rect 174262 11568 174268 11620
rect 174320 11608 174326 11620
rect 278958 11608 278964 11620
rect 174320 11580 278964 11608
rect 174320 11568 174326 11580
rect 278958 11568 278964 11580
rect 279016 11568 279022 11620
rect 177850 11500 177856 11552
rect 177908 11540 177914 11552
rect 279050 11540 279056 11552
rect 177908 11512 279056 11540
rect 177908 11500 177914 11512
rect 279050 11500 279056 11512
rect 279108 11500 279114 11552
rect 181438 11432 181444 11484
rect 181496 11472 181502 11484
rect 280522 11472 280528 11484
rect 181496 11444 280528 11472
rect 181496 11432 181502 11444
rect 280522 11432 280528 11444
rect 280580 11432 280586 11484
rect 184934 11364 184940 11416
rect 184992 11404 184998 11416
rect 281810 11404 281816 11416
rect 184992 11376 281816 11404
rect 184992 11364 184998 11376
rect 281810 11364 281816 11376
rect 281868 11364 281874 11416
rect 205542 11296 205548 11348
rect 205600 11336 205606 11348
rect 285950 11336 285956 11348
rect 205600 11308 285956 11336
rect 205600 11296 205606 11308
rect 285950 11296 285956 11308
rect 286008 11296 286014 11348
rect 209038 11228 209044 11280
rect 209096 11268 209102 11280
rect 287422 11268 287428 11280
rect 209096 11240 287428 11268
rect 209096 11228 209102 11240
rect 287422 11228 287428 11240
rect 287480 11228 287486 11280
rect 212166 11160 212172 11212
rect 212224 11200 212230 11212
rect 288710 11200 288716 11212
rect 212224 11172 288716 11200
rect 212224 11160 212230 11172
rect 288710 11160 288716 11172
rect 288768 11160 288774 11212
rect 215662 11092 215668 11144
rect 215720 11132 215726 11144
rect 288618 11132 288624 11144
rect 215720 11104 288624 11132
rect 215720 11092 215726 11104
rect 288618 11092 288624 11104
rect 288676 11092 288682 11144
rect 91002 10956 91008 11008
rect 91060 10996 91066 11008
rect 256878 10996 256884 11008
rect 91060 10968 256884 10996
rect 91060 10956 91066 10968
rect 256878 10956 256884 10968
rect 256936 10956 256942 11008
rect 357066 10956 357072 11008
rect 357124 10996 357130 11008
rect 480530 10996 480536 11008
rect 357124 10968 480536 10996
rect 357124 10956 357130 10968
rect 480530 10956 480536 10968
rect 480588 10956 480594 11008
rect 86678 10888 86684 10940
rect 86736 10928 86742 10940
rect 256786 10928 256792 10940
rect 86736 10900 256792 10928
rect 86736 10888 86742 10900
rect 256786 10888 256792 10900
rect 256844 10888 256850 10940
rect 357342 10888 357348 10940
rect 357400 10928 357406 10940
rect 481634 10928 481640 10940
rect 357400 10900 481640 10928
rect 357400 10888 357406 10900
rect 481634 10888 481640 10900
rect 481692 10888 481698 10940
rect 84102 10820 84108 10872
rect 84160 10860 84166 10872
rect 255590 10860 255596 10872
rect 84160 10832 255596 10860
rect 84160 10820 84166 10832
rect 255590 10820 255596 10832
rect 255648 10820 255654 10872
rect 357250 10820 357256 10872
rect 357308 10860 357314 10872
rect 481726 10860 481732 10872
rect 357308 10832 481732 10860
rect 357308 10820 357314 10832
rect 481726 10820 481732 10832
rect 481784 10820 481790 10872
rect 74442 10752 74448 10804
rect 74500 10792 74506 10804
rect 252738 10792 252744 10804
rect 74500 10764 252744 10792
rect 74500 10752 74506 10764
rect 252738 10752 252744 10764
rect 252796 10752 252802 10804
rect 358722 10752 358728 10804
rect 358780 10792 358786 10804
rect 484762 10792 484768 10804
rect 358780 10764 484768 10792
rect 358780 10752 358786 10764
rect 484762 10752 484768 10764
rect 484820 10752 484826 10804
rect 70302 10684 70308 10736
rect 70360 10724 70366 10736
rect 252830 10724 252836 10736
rect 70360 10696 252836 10724
rect 70360 10684 70366 10696
rect 252830 10684 252836 10696
rect 252888 10684 252894 10736
rect 357158 10684 357164 10736
rect 357216 10724 357222 10736
rect 484026 10724 484032 10736
rect 357216 10696 484032 10724
rect 357216 10684 357222 10696
rect 484026 10684 484032 10696
rect 484084 10684 484090 10736
rect 67542 10616 67548 10668
rect 67600 10656 67606 10668
rect 251450 10656 251456 10668
rect 67600 10628 251456 10656
rect 67600 10616 67606 10628
rect 251450 10616 251456 10628
rect 251508 10616 251514 10668
rect 358446 10616 358452 10668
rect 358504 10656 358510 10668
rect 486418 10656 486424 10668
rect 358504 10628 486424 10656
rect 358504 10616 358510 10628
rect 486418 10616 486424 10628
rect 486476 10616 486482 10668
rect 63218 10548 63224 10600
rect 63276 10588 63282 10600
rect 249886 10588 249892 10600
rect 63276 10560 249892 10588
rect 63276 10548 63282 10560
rect 249886 10548 249892 10560
rect 249944 10548 249950 10600
rect 358538 10548 358544 10600
rect 358596 10588 358602 10600
rect 487154 10588 487160 10600
rect 358596 10560 487160 10588
rect 358596 10548 358602 10560
rect 487154 10548 487160 10560
rect 487212 10548 487218 10600
rect 60642 10480 60648 10532
rect 60700 10520 60706 10532
rect 249978 10520 249984 10532
rect 60700 10492 249984 10520
rect 60700 10480 60706 10492
rect 249978 10480 249984 10492
rect 250036 10480 250042 10532
rect 358630 10480 358636 10532
rect 358688 10520 358694 10532
rect 488810 10520 488816 10532
rect 358688 10492 488816 10520
rect 358688 10480 358694 10492
rect 488810 10480 488816 10492
rect 488868 10480 488874 10532
rect 56502 10412 56508 10464
rect 56560 10452 56566 10464
rect 248414 10452 248420 10464
rect 56560 10424 248420 10452
rect 56560 10412 56566 10424
rect 248414 10412 248420 10424
rect 248472 10412 248478 10464
rect 359918 10412 359924 10464
rect 359976 10452 359982 10464
rect 490006 10452 490012 10464
rect 359976 10424 490012 10452
rect 359976 10412 359982 10424
rect 490006 10412 490012 10424
rect 490064 10412 490070 10464
rect 53650 10344 53656 10396
rect 53708 10384 53714 10396
rect 247310 10384 247316 10396
rect 53708 10356 247316 10384
rect 53708 10344 53714 10356
rect 247310 10344 247316 10356
rect 247368 10344 247374 10396
rect 359734 10344 359740 10396
rect 359792 10384 359798 10396
rect 489914 10384 489920 10396
rect 359792 10356 489920 10384
rect 359792 10344 359798 10356
rect 489914 10344 489920 10356
rect 489972 10344 489978 10396
rect 49602 10276 49608 10328
rect 49660 10316 49666 10328
rect 247402 10316 247408 10328
rect 49660 10288 247408 10316
rect 49660 10276 49666 10288
rect 247402 10276 247408 10288
rect 247460 10276 247466 10328
rect 359826 10276 359832 10328
rect 359884 10316 359890 10328
rect 493042 10316 493048 10328
rect 359884 10288 493048 10316
rect 359884 10276 359890 10288
rect 493042 10276 493048 10288
rect 493100 10276 493106 10328
rect 95050 10208 95056 10260
rect 95108 10248 95114 10260
rect 258166 10248 258172 10260
rect 95108 10220 258172 10248
rect 95108 10208 95114 10220
rect 258166 10208 258172 10220
rect 258224 10208 258230 10260
rect 355778 10208 355784 10260
rect 355836 10248 355842 10260
rect 476482 10248 476488 10260
rect 355836 10220 476488 10248
rect 355836 10208 355842 10220
rect 476482 10208 476488 10220
rect 476540 10208 476546 10260
rect 97902 10140 97908 10192
rect 97960 10180 97966 10192
rect 259546 10180 259552 10192
rect 97960 10152 259552 10180
rect 97960 10140 97966 10152
rect 259546 10140 259552 10152
rect 259604 10140 259610 10192
rect 355686 10140 355692 10192
rect 355744 10180 355750 10192
rect 473446 10180 473452 10192
rect 355744 10152 473452 10180
rect 355744 10140 355750 10152
rect 473446 10140 473452 10152
rect 473504 10140 473510 10192
rect 102042 10072 102048 10124
rect 102100 10112 102106 10124
rect 259822 10112 259828 10124
rect 102100 10084 259828 10112
rect 102100 10072 102106 10084
rect 259822 10072 259828 10084
rect 259880 10072 259886 10124
rect 355870 10072 355876 10124
rect 355928 10112 355934 10124
rect 473354 10112 473360 10124
rect 355928 10084 473360 10112
rect 355928 10072 355934 10084
rect 473354 10072 473360 10084
rect 473412 10072 473418 10124
rect 104526 10004 104532 10056
rect 104584 10044 104590 10056
rect 260926 10044 260932 10056
rect 104584 10016 260932 10044
rect 104584 10004 104590 10016
rect 260926 10004 260932 10016
rect 260984 10004 260990 10056
rect 334986 10004 334992 10056
rect 335044 10044 335050 10056
rect 395338 10044 395344 10056
rect 335044 10016 395344 10044
rect 335044 10004 335050 10016
rect 395338 10004 395344 10016
rect 395396 10004 395402 10056
rect 108942 9936 108948 9988
rect 109000 9976 109006 9988
rect 262306 9976 262312 9988
rect 109000 9948 262312 9976
rect 109000 9936 109006 9948
rect 262306 9936 262312 9948
rect 262364 9936 262370 9988
rect 334894 9936 334900 9988
rect 334952 9976 334958 9988
rect 392578 9976 392584 9988
rect 334952 9948 392584 9976
rect 334952 9936 334958 9948
rect 392578 9936 392584 9948
rect 392636 9936 392642 9988
rect 111610 9868 111616 9920
rect 111668 9908 111674 9920
rect 262398 9908 262404 9920
rect 111668 9880 262404 9908
rect 111668 9868 111674 9880
rect 262398 9868 262404 9880
rect 262456 9868 262462 9920
rect 335078 9868 335084 9920
rect 335136 9908 335142 9920
rect 391106 9908 391112 9920
rect 335136 9880 391112 9908
rect 335136 9868 335142 9880
rect 391106 9868 391112 9880
rect 391164 9868 391170 9920
rect 115842 9800 115848 9852
rect 115900 9840 115906 9852
rect 263686 9840 263692 9852
rect 115900 9812 263692 9840
rect 115900 9800 115906 9812
rect 263686 9800 263692 9812
rect 263744 9800 263750 9852
rect 333698 9800 333704 9852
rect 333756 9840 333762 9852
rect 389450 9840 389456 9852
rect 333756 9812 389456 9840
rect 333756 9800 333762 9812
rect 389450 9800 389456 9812
rect 389508 9800 389514 9852
rect 119798 9732 119804 9784
rect 119856 9772 119862 9784
rect 265250 9772 265256 9784
rect 119856 9744 265256 9772
rect 119856 9732 119862 9744
rect 265250 9732 265256 9744
rect 265308 9732 265314 9784
rect 333606 9732 333612 9784
rect 333664 9772 333670 9784
rect 387794 9772 387800 9784
rect 333664 9744 387800 9772
rect 333664 9732 333670 9744
rect 387794 9732 387800 9744
rect 387852 9732 387858 9784
rect 122742 9664 122748 9716
rect 122800 9704 122806 9716
rect 265066 9704 265072 9716
rect 122800 9676 265072 9704
rect 122800 9664 122806 9676
rect 265066 9664 265072 9676
rect 265124 9664 265130 9716
rect 332134 9664 332140 9716
rect 332192 9704 332198 9716
rect 384298 9704 384304 9716
rect 332192 9676 384304 9704
rect 332192 9664 332198 9676
rect 384298 9664 384304 9676
rect 384356 9664 384362 9716
rect 199102 9596 199108 9648
rect 199160 9636 199166 9648
rect 284570 9636 284576 9648
rect 199160 9608 284576 9636
rect 199160 9596 199166 9608
rect 284570 9596 284576 9608
rect 284628 9596 284634 9648
rect 343266 9596 343272 9648
rect 343324 9636 343330 9648
rect 428458 9636 428464 9648
rect 343324 9608 428464 9636
rect 343324 9596 343330 9608
rect 428458 9596 428464 9608
rect 428516 9596 428522 9648
rect 195606 9528 195612 9580
rect 195664 9568 195670 9580
rect 284662 9568 284668 9580
rect 195664 9540 284668 9568
rect 195664 9528 195670 9540
rect 284662 9528 284668 9540
rect 284720 9528 284726 9580
rect 344646 9528 344652 9580
rect 344704 9568 344710 9580
rect 432046 9568 432052 9580
rect 344704 9540 432052 9568
rect 344704 9528 344710 9540
rect 432046 9528 432052 9540
rect 432104 9528 432110 9580
rect 192018 9460 192024 9512
rect 192076 9500 192082 9512
rect 283282 9500 283288 9512
rect 192076 9472 283288 9500
rect 192076 9460 192082 9472
rect 283282 9460 283288 9472
rect 283340 9460 283346 9512
rect 346026 9460 346032 9512
rect 346084 9500 346090 9512
rect 435542 9500 435548 9512
rect 346084 9472 435548 9500
rect 346084 9460 346090 9472
rect 435542 9460 435548 9472
rect 435600 9460 435606 9512
rect 188522 9392 188528 9444
rect 188580 9432 188586 9444
rect 281718 9432 281724 9444
rect 188580 9404 281724 9432
rect 188580 9392 188586 9404
rect 281718 9392 281724 9404
rect 281776 9392 281782 9444
rect 346118 9392 346124 9444
rect 346176 9432 346182 9444
rect 439130 9432 439136 9444
rect 346176 9404 439136 9432
rect 346176 9392 346182 9404
rect 439130 9392 439136 9404
rect 439188 9392 439194 9444
rect 156598 9324 156604 9376
rect 156656 9364 156662 9376
rect 273622 9364 273628 9376
rect 156656 9336 273628 9364
rect 156656 9324 156662 9336
rect 273622 9324 273628 9336
rect 273680 9324 273686 9376
rect 347406 9324 347412 9376
rect 347464 9364 347470 9376
rect 442626 9364 442632 9376
rect 347464 9336 442632 9364
rect 347464 9324 347470 9336
rect 442626 9324 442632 9336
rect 442684 9324 442690 9376
rect 153010 9256 153016 9308
rect 153068 9296 153074 9308
rect 273530 9296 273536 9308
rect 153068 9268 273536 9296
rect 153068 9256 153074 9268
rect 273530 9256 273536 9268
rect 273588 9256 273594 9308
rect 348878 9256 348884 9308
rect 348936 9296 348942 9308
rect 446214 9296 446220 9308
rect 348936 9268 446220 9296
rect 348936 9256 348942 9268
rect 446214 9256 446220 9268
rect 446272 9256 446278 9308
rect 149514 9188 149520 9240
rect 149572 9228 149578 9240
rect 272058 9228 272064 9240
rect 149572 9200 272064 9228
rect 149572 9188 149578 9200
rect 272058 9188 272064 9200
rect 272116 9188 272122 9240
rect 348970 9188 348976 9240
rect 349028 9228 349034 9240
rect 449802 9228 449808 9240
rect 349028 9200 449808 9228
rect 349028 9188 349034 9200
rect 449802 9188 449808 9200
rect 449860 9188 449866 9240
rect 145926 9120 145932 9172
rect 145984 9160 145990 9172
rect 270770 9160 270776 9172
rect 145984 9132 270776 9160
rect 145984 9120 145990 9132
rect 270770 9120 270776 9132
rect 270828 9120 270834 9172
rect 350258 9120 350264 9172
rect 350316 9160 350322 9172
rect 453298 9160 453304 9172
rect 350316 9132 453304 9160
rect 350316 9120 350322 9132
rect 453298 9120 453304 9132
rect 453356 9120 453362 9172
rect 142430 9052 142436 9104
rect 142488 9092 142494 9104
rect 270678 9092 270684 9104
rect 142488 9064 270684 9092
rect 142488 9052 142494 9064
rect 270678 9052 270684 9064
rect 270736 9052 270742 9104
rect 351546 9052 351552 9104
rect 351604 9092 351610 9104
rect 456886 9092 456892 9104
rect 351604 9064 456892 9092
rect 351604 9052 351610 9064
rect 456886 9052 456892 9064
rect 456944 9052 456950 9104
rect 138842 8984 138848 9036
rect 138900 9024 138906 9036
rect 269206 9024 269212 9036
rect 138900 8996 269212 9024
rect 138900 8984 138906 8996
rect 269206 8984 269212 8996
rect 269264 8984 269270 9036
rect 351638 8984 351644 9036
rect 351696 9024 351702 9036
rect 460382 9024 460388 9036
rect 351696 8996 460388 9024
rect 351696 8984 351702 8996
rect 460382 8984 460388 8996
rect 460440 8984 460446 9036
rect 33594 8916 33600 8968
rect 33652 8956 33658 8968
rect 242986 8956 242992 8968
rect 33652 8928 242992 8956
rect 33652 8916 33658 8928
rect 242986 8916 242992 8928
rect 243044 8916 243050 8968
rect 248782 8916 248788 8968
rect 248840 8956 248846 8968
rect 296898 8956 296904 8968
rect 248840 8928 296904 8956
rect 248840 8916 248846 8928
rect 296898 8916 296904 8928
rect 296956 8916 296962 8968
rect 352834 8916 352840 8968
rect 352892 8956 352898 8968
rect 463970 8956 463976 8968
rect 352892 8928 463976 8956
rect 352892 8916 352898 8928
rect 463970 8916 463976 8928
rect 464028 8916 464034 8968
rect 202690 8848 202696 8900
rect 202748 8888 202754 8900
rect 285858 8888 285864 8900
rect 202748 8860 285864 8888
rect 202748 8848 202754 8860
rect 285858 8848 285864 8860
rect 285916 8848 285922 8900
rect 343358 8848 343364 8900
rect 343416 8888 343422 8900
rect 424962 8888 424968 8900
rect 343416 8860 424968 8888
rect 343416 8848 343422 8860
rect 424962 8848 424968 8860
rect 425020 8848 425026 8900
rect 206186 8780 206192 8832
rect 206244 8820 206250 8832
rect 287238 8820 287244 8832
rect 206244 8792 287244 8820
rect 206244 8780 206250 8792
rect 287238 8780 287244 8792
rect 287296 8780 287302 8832
rect 341978 8780 341984 8832
rect 342036 8820 342042 8832
rect 421374 8820 421380 8832
rect 342036 8792 421380 8820
rect 342036 8780 342042 8792
rect 421374 8780 421380 8792
rect 421432 8780 421438 8832
rect 209774 8712 209780 8764
rect 209832 8752 209838 8764
rect 287330 8752 287336 8764
rect 209832 8724 287336 8752
rect 209832 8712 209838 8724
rect 287330 8712 287336 8724
rect 287388 8712 287394 8764
rect 340598 8712 340604 8764
rect 340656 8752 340662 8764
rect 417878 8752 417884 8764
rect 340656 8724 417884 8752
rect 340656 8712 340662 8724
rect 417878 8712 417884 8724
rect 417936 8712 417942 8764
rect 213362 8644 213368 8696
rect 213420 8684 213426 8696
rect 288526 8684 288532 8696
rect 213420 8656 288532 8684
rect 213420 8644 213426 8656
rect 288526 8644 288532 8656
rect 288584 8644 288590 8696
rect 340690 8644 340696 8696
rect 340748 8684 340754 8696
rect 414290 8684 414296 8696
rect 340748 8656 414296 8684
rect 340748 8644 340754 8656
rect 414290 8644 414296 8656
rect 414348 8644 414354 8696
rect 216858 8576 216864 8628
rect 216916 8616 216922 8628
rect 289998 8616 290004 8628
rect 216916 8588 290004 8616
rect 216916 8576 216922 8588
rect 289998 8576 290004 8588
rect 290056 8576 290062 8628
rect 339126 8576 339132 8628
rect 339184 8616 339190 8628
rect 410794 8616 410800 8628
rect 339184 8588 410800 8616
rect 339184 8576 339190 8588
rect 410794 8576 410800 8588
rect 410852 8576 410858 8628
rect 220446 8508 220452 8560
rect 220504 8548 220510 8560
rect 289906 8548 289912 8560
rect 220504 8520 289912 8548
rect 220504 8508 220510 8520
rect 289906 8508 289912 8520
rect 289964 8508 289970 8560
rect 337746 8508 337752 8560
rect 337804 8548 337810 8560
rect 407206 8548 407212 8560
rect 337804 8520 407212 8548
rect 337804 8508 337810 8520
rect 407206 8508 407212 8520
rect 407264 8508 407270 8560
rect 223942 8440 223948 8492
rect 224000 8480 224006 8492
rect 291562 8480 291568 8492
rect 224000 8452 291568 8480
rect 224000 8440 224006 8452
rect 291562 8440 291568 8452
rect 291620 8440 291626 8492
rect 337838 8440 337844 8492
rect 337896 8480 337902 8492
rect 403526 8480 403532 8492
rect 337896 8452 403532 8480
rect 337896 8440 337902 8452
rect 403526 8440 403532 8452
rect 403584 8440 403590 8492
rect 227530 8372 227536 8424
rect 227588 8412 227594 8424
rect 291470 8412 291476 8424
rect 227588 8384 291476 8412
rect 227588 8372 227594 8384
rect 291470 8372 291476 8384
rect 291528 8372 291534 8424
rect 336366 8372 336372 8424
rect 336424 8412 336430 8424
rect 400122 8412 400128 8424
rect 336424 8384 400128 8412
rect 336424 8372 336430 8384
rect 400122 8372 400128 8384
rect 400180 8372 400186 8424
rect 231026 8304 231032 8356
rect 231084 8344 231090 8356
rect 292850 8344 292856 8356
rect 231084 8316 292856 8344
rect 231084 8304 231090 8316
rect 292850 8304 292856 8316
rect 292908 8304 292914 8356
rect 335170 8304 335176 8356
rect 335228 8344 335234 8356
rect 396534 8344 396540 8356
rect 335228 8316 396540 8344
rect 335228 8304 335234 8316
rect 396534 8304 396540 8316
rect 396592 8304 396598 8356
rect 151814 8236 151820 8288
rect 151872 8276 151878 8288
rect 273346 8276 273352 8288
rect 151872 8248 273352 8276
rect 151872 8236 151878 8248
rect 273346 8236 273352 8248
rect 273404 8236 273410 8288
rect 366818 8236 366824 8288
rect 366876 8276 366882 8288
rect 520734 8276 520740 8288
rect 366876 8248 520740 8276
rect 366876 8236 366882 8248
rect 520734 8236 520740 8248
rect 520792 8236 520798 8288
rect 148318 8168 148324 8220
rect 148376 8208 148382 8220
rect 271966 8208 271972 8220
rect 148376 8180 271972 8208
rect 148376 8168 148382 8180
rect 271966 8168 271972 8180
rect 272024 8168 272030 8220
rect 368198 8168 368204 8220
rect 368256 8208 368262 8220
rect 524230 8208 524236 8220
rect 368256 8180 524236 8208
rect 368256 8168 368262 8180
rect 524230 8168 524236 8180
rect 524288 8168 524294 8220
rect 144730 8100 144736 8152
rect 144788 8140 144794 8152
rect 270586 8140 270592 8152
rect 144788 8112 270592 8140
rect 144788 8100 144794 8112
rect 270586 8100 270592 8112
rect 270644 8100 270650 8152
rect 369486 8100 369492 8152
rect 369544 8140 369550 8152
rect 527818 8140 527824 8152
rect 369544 8112 527824 8140
rect 369544 8100 369550 8112
rect 527818 8100 527824 8112
rect 527876 8100 527882 8152
rect 141234 8032 141240 8084
rect 141292 8072 141298 8084
rect 270494 8072 270500 8084
rect 141292 8044 270500 8072
rect 141292 8032 141298 8044
rect 270494 8032 270500 8044
rect 270552 8032 270558 8084
rect 369578 8032 369584 8084
rect 369636 8072 369642 8084
rect 531314 8072 531320 8084
rect 369636 8044 531320 8072
rect 369636 8032 369642 8044
rect 531314 8032 531320 8044
rect 531372 8032 531378 8084
rect 137646 7964 137652 8016
rect 137704 8004 137710 8016
rect 269114 8004 269120 8016
rect 137704 7976 269120 8004
rect 137704 7964 137710 7976
rect 269114 7964 269120 7976
rect 269172 7964 269178 8016
rect 370866 7964 370872 8016
rect 370924 8004 370930 8016
rect 534902 8004 534908 8016
rect 370924 7976 534908 8004
rect 370924 7964 370930 7976
rect 534902 7964 534908 7976
rect 534960 7964 534966 8016
rect 134150 7896 134156 7948
rect 134208 7936 134214 7948
rect 267918 7936 267924 7948
rect 134208 7908 267924 7936
rect 134208 7896 134214 7908
rect 267918 7896 267924 7908
rect 267976 7896 267982 7948
rect 370958 7896 370964 7948
rect 371016 7936 371022 7948
rect 538398 7936 538404 7948
rect 371016 7908 538404 7936
rect 371016 7896 371022 7908
rect 538398 7896 538404 7908
rect 538456 7896 538462 7948
rect 128170 7828 128176 7880
rect 128228 7868 128234 7880
rect 266538 7868 266544 7880
rect 128228 7840 266544 7868
rect 128228 7828 128234 7840
rect 266538 7828 266544 7840
rect 266596 7828 266602 7880
rect 372430 7828 372436 7880
rect 372488 7868 372494 7880
rect 541986 7868 541992 7880
rect 372488 7840 541992 7868
rect 372488 7828 372494 7840
rect 541986 7828 541992 7840
rect 542044 7828 542050 7880
rect 76190 7760 76196 7812
rect 76248 7800 76254 7812
rect 249705 7803 249763 7809
rect 249705 7800 249717 7803
rect 76248 7772 249717 7800
rect 76248 7760 76254 7772
rect 249705 7769 249717 7772
rect 249751 7769 249763 7803
rect 252646 7800 252652 7812
rect 249705 7763 249763 7769
rect 249812 7772 252652 7800
rect 72602 7692 72608 7744
rect 72660 7732 72666 7744
rect 249812 7732 249840 7772
rect 252646 7760 252652 7772
rect 252704 7760 252710 7812
rect 261754 7760 261760 7812
rect 261812 7800 261818 7812
rect 301038 7800 301044 7812
rect 261812 7772 301044 7800
rect 261812 7760 261818 7772
rect 301038 7760 301044 7772
rect 301096 7760 301102 7812
rect 373626 7760 373632 7812
rect 373684 7800 373690 7812
rect 545482 7800 545488 7812
rect 373684 7772 545488 7800
rect 373684 7760 373690 7772
rect 545482 7760 545488 7772
rect 545540 7760 545546 7812
rect 251358 7732 251364 7744
rect 72660 7704 249840 7732
rect 249996 7704 251364 7732
rect 72660 7692 72666 7704
rect 69106 7624 69112 7676
rect 69164 7664 69170 7676
rect 249889 7667 249947 7673
rect 249889 7664 249901 7667
rect 69164 7636 249901 7664
rect 69164 7624 69170 7636
rect 249889 7633 249901 7636
rect 249935 7633 249947 7667
rect 249889 7627 249947 7633
rect 65518 7556 65524 7608
rect 65576 7596 65582 7608
rect 249996 7596 250024 7704
rect 251358 7692 251364 7704
rect 251416 7692 251422 7744
rect 258258 7692 258264 7744
rect 258316 7732 258322 7744
rect 299566 7732 299572 7744
rect 258316 7704 299572 7732
rect 258316 7692 258322 7704
rect 299566 7692 299572 7704
rect 299624 7692 299630 7744
rect 373718 7692 373724 7744
rect 373776 7732 373782 7744
rect 549070 7732 549076 7744
rect 373776 7704 549076 7732
rect 373776 7692 373782 7704
rect 549070 7692 549076 7704
rect 549128 7692 549134 7744
rect 250073 7667 250131 7673
rect 250073 7633 250085 7667
rect 250119 7664 250131 7667
rect 251266 7664 251272 7676
rect 250119 7636 251272 7664
rect 250119 7633 250131 7636
rect 250073 7627 250131 7633
rect 251266 7624 251272 7636
rect 251324 7624 251330 7676
rect 254670 7624 254676 7676
rect 254728 7664 254734 7676
rect 298278 7664 298284 7676
rect 254728 7636 298284 7664
rect 254728 7624 254734 7636
rect 298278 7624 298284 7636
rect 298336 7624 298342 7676
rect 374914 7624 374920 7676
rect 374972 7664 374978 7676
rect 552658 7664 552664 7676
rect 374972 7636 552664 7664
rect 374972 7624 374978 7636
rect 552658 7624 552664 7636
rect 552716 7624 552722 7676
rect 65576 7568 250024 7596
rect 65576 7556 65582 7568
rect 251174 7556 251180 7608
rect 251232 7596 251238 7608
rect 298370 7596 298376 7608
rect 251232 7568 298376 7596
rect 251232 7556 251238 7568
rect 298370 7556 298376 7568
rect 298428 7556 298434 7608
rect 376478 7556 376484 7608
rect 376536 7596 376542 7608
rect 556154 7596 556160 7608
rect 376536 7568 556160 7596
rect 376536 7556 376542 7568
rect 556154 7556 556160 7568
rect 556212 7556 556218 7608
rect 155402 7488 155408 7540
rect 155460 7528 155466 7540
rect 273438 7528 273444 7540
rect 155460 7500 273444 7528
rect 155460 7488 155466 7500
rect 273438 7488 273444 7500
rect 273496 7488 273502 7540
rect 366910 7488 366916 7540
rect 366968 7528 366974 7540
rect 517146 7528 517152 7540
rect 366968 7500 517152 7528
rect 366968 7488 366974 7500
rect 517146 7488 517152 7500
rect 517204 7488 517210 7540
rect 158898 7420 158904 7472
rect 158956 7460 158962 7472
rect 274726 7460 274732 7472
rect 158956 7432 274732 7460
rect 158956 7420 158962 7432
rect 274726 7420 274732 7432
rect 274784 7420 274790 7472
rect 365438 7420 365444 7472
rect 365496 7460 365502 7472
rect 513558 7460 513564 7472
rect 365496 7432 513564 7460
rect 365496 7420 365502 7432
rect 513558 7420 513564 7432
rect 513616 7420 513622 7472
rect 163682 7352 163688 7404
rect 163740 7392 163746 7404
rect 276290 7392 276296 7404
rect 163740 7364 276296 7392
rect 163740 7352 163746 7364
rect 276290 7352 276296 7364
rect 276348 7352 276354 7404
rect 364058 7352 364064 7404
rect 364116 7392 364122 7404
rect 510062 7392 510068 7404
rect 364116 7364 510068 7392
rect 364116 7352 364122 7364
rect 510062 7352 510068 7364
rect 510120 7352 510126 7404
rect 167178 7284 167184 7336
rect 167236 7324 167242 7336
rect 276198 7324 276204 7336
rect 167236 7296 276204 7324
rect 167236 7284 167242 7296
rect 276198 7284 276204 7296
rect 276256 7284 276262 7336
rect 364150 7284 364156 7336
rect 364208 7324 364214 7336
rect 506474 7324 506480 7336
rect 364208 7296 506480 7324
rect 364208 7284 364214 7296
rect 506474 7284 506480 7296
rect 506532 7284 506538 7336
rect 170766 7216 170772 7268
rect 170824 7256 170830 7268
rect 277578 7256 277584 7268
rect 170824 7228 277584 7256
rect 170824 7216 170830 7228
rect 277578 7216 277584 7228
rect 277636 7216 277642 7268
rect 362678 7216 362684 7268
rect 362736 7256 362742 7268
rect 502978 7256 502984 7268
rect 362736 7228 502984 7256
rect 362736 7216 362742 7228
rect 502978 7216 502984 7228
rect 503036 7216 503042 7268
rect 222746 7148 222752 7200
rect 222804 7188 222810 7200
rect 291378 7188 291384 7200
rect 222804 7160 291384 7188
rect 222804 7148 222810 7160
rect 291378 7148 291384 7160
rect 291436 7148 291442 7200
rect 361390 7148 361396 7200
rect 361448 7188 361454 7200
rect 499390 7188 499396 7200
rect 361448 7160 499396 7188
rect 361448 7148 361454 7160
rect 499390 7148 499396 7160
rect 499448 7148 499454 7200
rect 229830 7080 229836 7132
rect 229888 7120 229894 7132
rect 292758 7120 292764 7132
rect 229888 7092 292764 7120
rect 229888 7080 229894 7092
rect 292758 7080 292764 7092
rect 292816 7080 292822 7132
rect 361298 7080 361304 7132
rect 361356 7120 361362 7132
rect 495894 7120 495900 7132
rect 361356 7092 495900 7120
rect 361356 7080 361362 7092
rect 495894 7080 495900 7092
rect 495952 7080 495958 7132
rect 233418 7012 233424 7064
rect 233476 7052 233482 7064
rect 294322 7052 294328 7064
rect 233476 7024 294328 7052
rect 233476 7012 233482 7024
rect 294322 7012 294328 7024
rect 294380 7012 294386 7064
rect 360102 7012 360108 7064
rect 360160 7052 360166 7064
rect 492306 7052 492312 7064
rect 360160 7024 492312 7052
rect 360160 7012 360166 7024
rect 492306 7012 492312 7024
rect 492364 7012 492370 7064
rect 219250 6944 219256 6996
rect 219308 6984 219314 6996
rect 246298 6984 246304 6996
rect 219308 6956 246304 6984
rect 219308 6944 219314 6956
rect 246298 6944 246304 6956
rect 246356 6944 246362 6996
rect 247586 6944 247592 6996
rect 247644 6984 247650 6996
rect 296806 6984 296812 6996
rect 247644 6956 296812 6984
rect 247644 6944 247650 6956
rect 296806 6944 296812 6956
rect 296864 6944 296870 6996
rect 332226 6944 332232 6996
rect 332284 6984 332290 6996
rect 385954 6984 385960 6996
rect 332284 6956 385960 6984
rect 332284 6944 332290 6956
rect 385954 6944 385960 6956
rect 386012 6944 386018 6996
rect 249705 6919 249763 6925
rect 249705 6885 249717 6919
rect 249751 6916 249763 6919
rect 254026 6916 254032 6928
rect 249751 6888 254032 6916
rect 249751 6885 249763 6888
rect 249705 6879 249763 6885
rect 254026 6876 254032 6888
rect 254084 6876 254090 6928
rect 173158 6808 173164 6860
rect 173216 6848 173222 6860
rect 277670 6848 277676 6860
rect 173216 6820 277676 6848
rect 173216 6808 173222 6820
rect 277670 6808 277676 6820
rect 277728 6808 277734 6860
rect 332318 6808 332324 6860
rect 332376 6848 332382 6860
rect 382366 6848 382372 6860
rect 332376 6820 382372 6848
rect 332376 6808 332382 6820
rect 382366 6808 382372 6820
rect 382424 6808 382430 6860
rect 393958 6808 393964 6860
rect 394016 6848 394022 6860
rect 580166 6848 580172 6860
rect 394016 6820 580172 6848
rect 394016 6808 394022 6820
rect 580166 6808 580172 6820
rect 580224 6808 580230 6860
rect 169570 6740 169576 6792
rect 169628 6780 169634 6792
rect 277486 6780 277492 6792
rect 169628 6752 277492 6780
rect 169628 6740 169634 6752
rect 277486 6740 277492 6752
rect 277544 6740 277550 6792
rect 344738 6740 344744 6792
rect 344796 6780 344802 6792
rect 430850 6780 430856 6792
rect 344796 6752 430856 6780
rect 344796 6740 344802 6752
rect 430850 6740 430856 6752
rect 430908 6740 430914 6792
rect 166074 6672 166080 6724
rect 166132 6712 166138 6724
rect 276106 6712 276112 6724
rect 166132 6684 276112 6712
rect 166132 6672 166138 6684
rect 276106 6672 276112 6684
rect 276164 6672 276170 6724
rect 344830 6672 344836 6724
rect 344888 6712 344894 6724
rect 434438 6712 434444 6724
rect 344888 6684 434444 6712
rect 344888 6672 344894 6684
rect 434438 6672 434444 6684
rect 434496 6672 434502 6724
rect 3418 6604 3424 6656
rect 3476 6644 3482 6656
rect 7558 6644 7564 6656
rect 3476 6616 7564 6644
rect 3476 6604 3482 6616
rect 7558 6604 7564 6616
rect 7616 6604 7622 6656
rect 162486 6604 162492 6656
rect 162544 6644 162550 6656
rect 276014 6644 276020 6656
rect 162544 6616 276020 6644
rect 162544 6604 162550 6616
rect 276014 6604 276020 6616
rect 276072 6604 276078 6656
rect 346210 6604 346216 6656
rect 346268 6644 346274 6656
rect 437934 6644 437940 6656
rect 346268 6616 437940 6644
rect 346268 6604 346274 6616
rect 437934 6604 437940 6616
rect 437992 6604 437998 6656
rect 157794 6536 157800 6588
rect 157852 6576 157858 6588
rect 274634 6576 274640 6588
rect 157852 6548 274640 6576
rect 157852 6536 157858 6548
rect 274634 6536 274640 6548
rect 274692 6536 274698 6588
rect 347498 6536 347504 6588
rect 347556 6576 347562 6588
rect 441522 6576 441528 6588
rect 347556 6548 441528 6576
rect 347556 6536 347562 6548
rect 441522 6536 441528 6548
rect 441580 6536 441586 6588
rect 154206 6468 154212 6520
rect 154264 6508 154270 6520
rect 273254 6508 273260 6520
rect 154264 6480 273260 6508
rect 154264 6468 154270 6480
rect 273254 6468 273260 6480
rect 273312 6468 273318 6520
rect 347590 6468 347596 6520
rect 347648 6508 347654 6520
rect 445018 6508 445024 6520
rect 347648 6480 445024 6508
rect 347648 6468 347654 6480
rect 445018 6468 445024 6480
rect 445076 6468 445082 6520
rect 150618 6400 150624 6452
rect 150676 6440 150682 6452
rect 271874 6440 271880 6452
rect 150676 6412 271880 6440
rect 150676 6400 150682 6412
rect 271874 6400 271880 6412
rect 271932 6400 271938 6452
rect 349062 6400 349068 6452
rect 349120 6440 349126 6452
rect 448606 6440 448612 6452
rect 349120 6412 448612 6440
rect 349120 6400 349126 6412
rect 448606 6400 448612 6412
rect 448664 6400 448670 6452
rect 130562 6332 130568 6384
rect 130620 6372 130626 6384
rect 267826 6372 267832 6384
rect 130620 6344 267832 6372
rect 130620 6332 130626 6344
rect 267826 6332 267832 6344
rect 267884 6332 267890 6384
rect 350442 6332 350448 6384
rect 350500 6372 350506 6384
rect 452102 6372 452108 6384
rect 350500 6344 452108 6372
rect 350500 6332 350506 6344
rect 452102 6332 452108 6344
rect 452160 6332 452166 6384
rect 126974 6264 126980 6316
rect 127032 6304 127038 6316
rect 266446 6304 266452 6316
rect 127032 6276 266452 6304
rect 127032 6264 127038 6276
rect 266446 6264 266452 6276
rect 266504 6264 266510 6316
rect 350350 6264 350356 6316
rect 350408 6304 350414 6316
rect 455690 6304 455696 6316
rect 350408 6276 455696 6304
rect 350408 6264 350414 6276
rect 455690 6264 455696 6276
rect 455748 6264 455754 6316
rect 61930 6196 61936 6248
rect 61988 6236 61994 6248
rect 250070 6236 250076 6248
rect 61988 6208 250076 6236
rect 61988 6196 61994 6208
rect 250070 6196 250076 6208
rect 250128 6196 250134 6248
rect 351730 6196 351736 6248
rect 351788 6236 351794 6248
rect 459186 6236 459192 6248
rect 351788 6208 459192 6236
rect 351788 6196 351794 6208
rect 459186 6196 459192 6208
rect 459244 6196 459250 6248
rect 4062 6128 4068 6180
rect 4120 6168 4126 6180
rect 234890 6168 234896 6180
rect 4120 6140 234896 6168
rect 4120 6128 4126 6140
rect 234890 6128 234896 6140
rect 234948 6128 234954 6180
rect 238110 6128 238116 6180
rect 238168 6168 238174 6180
rect 294230 6168 294236 6180
rect 238168 6140 294236 6168
rect 238168 6128 238174 6140
rect 294230 6128 294236 6140
rect 294288 6128 294294 6180
rect 353110 6128 353116 6180
rect 353168 6168 353174 6180
rect 462774 6168 462780 6180
rect 353168 6140 462780 6168
rect 353168 6128 353174 6140
rect 462774 6128 462780 6140
rect 462832 6128 462838 6180
rect 176654 6060 176660 6112
rect 176712 6100 176718 6112
rect 278866 6100 278872 6112
rect 176712 6072 278872 6100
rect 176712 6060 176718 6072
rect 278866 6060 278872 6072
rect 278924 6060 278930 6112
rect 343450 6060 343456 6112
rect 343508 6100 343514 6112
rect 427262 6100 427268 6112
rect 343508 6072 427268 6100
rect 343508 6060 343514 6072
rect 427262 6060 427268 6072
rect 427320 6060 427326 6112
rect 180242 5992 180248 6044
rect 180300 6032 180306 6044
rect 280338 6032 280344 6044
rect 180300 6004 280344 6032
rect 180300 5992 180306 6004
rect 280338 5992 280344 6004
rect 280396 5992 280402 6044
rect 342070 5992 342076 6044
rect 342128 6032 342134 6044
rect 423766 6032 423772 6044
rect 342128 6004 423772 6032
rect 342128 5992 342134 6004
rect 423766 5992 423772 6004
rect 423824 5992 423830 6044
rect 183738 5924 183744 5976
rect 183796 5964 183802 5976
rect 280430 5964 280436 5976
rect 183796 5936 280436 5964
rect 183796 5924 183802 5936
rect 280430 5924 280436 5936
rect 280488 5924 280494 5976
rect 342162 5924 342168 5976
rect 342220 5964 342226 5976
rect 420178 5964 420184 5976
rect 342220 5936 420184 5964
rect 342220 5924 342226 5936
rect 420178 5924 420184 5936
rect 420236 5924 420242 5976
rect 187326 5856 187332 5908
rect 187384 5896 187390 5908
rect 281626 5896 281632 5908
rect 187384 5868 281632 5896
rect 187384 5856 187390 5868
rect 281626 5856 281632 5868
rect 281684 5856 281690 5908
rect 340782 5856 340788 5908
rect 340840 5896 340846 5908
rect 416682 5896 416688 5908
rect 340840 5868 416688 5896
rect 340840 5856 340846 5868
rect 416682 5856 416688 5868
rect 416740 5856 416746 5908
rect 190822 5788 190828 5840
rect 190880 5828 190886 5840
rect 283190 5828 283196 5840
rect 190880 5800 283196 5828
rect 190880 5788 190886 5800
rect 283190 5788 283196 5800
rect 283248 5788 283254 5840
rect 339310 5788 339316 5840
rect 339368 5828 339374 5840
rect 413094 5828 413100 5840
rect 339368 5800 413100 5828
rect 339368 5788 339374 5800
rect 413094 5788 413100 5800
rect 413152 5788 413158 5840
rect 194410 5720 194416 5772
rect 194468 5760 194474 5772
rect 283098 5760 283104 5772
rect 194468 5732 283104 5760
rect 194468 5720 194474 5732
rect 283098 5720 283104 5732
rect 283156 5720 283162 5772
rect 339218 5720 339224 5772
rect 339276 5760 339282 5772
rect 409598 5760 409604 5772
rect 339276 5732 409604 5760
rect 339276 5720 339282 5732
rect 409598 5720 409604 5732
rect 409656 5720 409662 5772
rect 197906 5652 197912 5704
rect 197964 5692 197970 5704
rect 284478 5692 284484 5704
rect 197964 5664 284484 5692
rect 197964 5652 197970 5664
rect 284478 5652 284484 5664
rect 284536 5652 284542 5704
rect 338022 5652 338028 5704
rect 338080 5692 338086 5704
rect 406010 5692 406016 5704
rect 338080 5664 406016 5692
rect 338080 5652 338086 5664
rect 406010 5652 406016 5664
rect 406068 5652 406074 5704
rect 201494 5584 201500 5636
rect 201552 5624 201558 5636
rect 285766 5624 285772 5636
rect 201552 5596 285772 5624
rect 201552 5584 201558 5596
rect 285766 5584 285772 5596
rect 285824 5584 285830 5636
rect 337930 5584 337936 5636
rect 337988 5624 337994 5636
rect 402514 5624 402520 5636
rect 337988 5596 402520 5624
rect 337988 5584 337994 5596
rect 402514 5584 402520 5596
rect 402572 5584 402578 5636
rect 226334 5516 226340 5568
rect 226392 5556 226398 5568
rect 291286 5556 291292 5568
rect 226392 5528 291292 5556
rect 226392 5516 226398 5528
rect 291286 5516 291292 5528
rect 291344 5516 291350 5568
rect 336458 5516 336464 5568
rect 336516 5556 336522 5568
rect 398926 5556 398932 5568
rect 336516 5528 398932 5556
rect 336516 5516 336522 5528
rect 398926 5516 398932 5528
rect 398984 5516 398990 5568
rect 203886 5448 203892 5500
rect 203944 5488 203950 5500
rect 285674 5488 285680 5500
rect 203944 5460 285680 5488
rect 203944 5448 203950 5460
rect 285674 5448 285680 5460
rect 285732 5448 285738 5500
rect 326706 5448 326712 5500
rect 326764 5488 326770 5500
rect 359918 5488 359924 5500
rect 326764 5460 359924 5488
rect 326764 5448 326770 5460
rect 359918 5448 359924 5460
rect 359976 5448 359982 5500
rect 368382 5448 368388 5500
rect 368440 5488 368446 5500
rect 526622 5488 526628 5500
rect 368440 5460 526628 5488
rect 368440 5448 368446 5460
rect 526622 5448 526628 5460
rect 526680 5448 526686 5500
rect 200298 5380 200304 5432
rect 200356 5420 200362 5432
rect 284386 5420 284392 5432
rect 200356 5392 284392 5420
rect 200356 5380 200362 5392
rect 284386 5380 284392 5392
rect 284444 5380 284450 5432
rect 326798 5380 326804 5432
rect 326856 5420 326862 5432
rect 361114 5420 361120 5432
rect 326856 5392 361120 5420
rect 326856 5380 326862 5392
rect 361114 5380 361120 5392
rect 361172 5380 361178 5432
rect 369670 5380 369676 5432
rect 369728 5420 369734 5432
rect 530118 5420 530124 5432
rect 369728 5392 530124 5420
rect 369728 5380 369734 5392
rect 530118 5380 530124 5392
rect 530176 5380 530182 5432
rect 123478 5312 123484 5364
rect 123536 5352 123542 5364
rect 191098 5352 191104 5364
rect 123536 5324 191104 5352
rect 123536 5312 123542 5324
rect 191098 5312 191104 5324
rect 191156 5312 191162 5364
rect 193214 5312 193220 5364
rect 193272 5352 193278 5364
rect 193272 5324 193996 5352
rect 193272 5312 193278 5324
rect 124674 5244 124680 5296
rect 124732 5284 124738 5296
rect 193858 5284 193864 5296
rect 124732 5256 193864 5284
rect 124732 5244 124738 5256
rect 193858 5244 193864 5256
rect 193916 5244 193922 5296
rect 193968 5284 193996 5324
rect 196802 5312 196808 5364
rect 196860 5352 196866 5364
rect 284294 5352 284300 5364
rect 196860 5324 284300 5352
rect 196860 5312 196866 5324
rect 284294 5312 284300 5324
rect 284352 5312 284358 5364
rect 328086 5312 328092 5364
rect 328144 5352 328150 5364
rect 364610 5352 364616 5364
rect 328144 5324 364616 5352
rect 328144 5312 328150 5324
rect 364610 5312 364616 5324
rect 364668 5312 364674 5364
rect 371050 5312 371056 5364
rect 371108 5352 371114 5364
rect 533706 5352 533712 5364
rect 371108 5324 533712 5352
rect 371108 5312 371114 5324
rect 533706 5312 533712 5324
rect 533764 5312 533770 5364
rect 283006 5284 283012 5296
rect 193968 5256 283012 5284
rect 283006 5244 283012 5256
rect 283064 5244 283070 5296
rect 326614 5244 326620 5296
rect 326672 5284 326678 5296
rect 363506 5284 363512 5296
rect 326672 5256 363512 5284
rect 326672 5244 326678 5256
rect 363506 5244 363512 5256
rect 363564 5244 363570 5296
rect 371142 5244 371148 5296
rect 371200 5284 371206 5296
rect 537202 5284 537208 5296
rect 371200 5256 537208 5284
rect 371200 5244 371206 5256
rect 537202 5244 537208 5256
rect 537260 5244 537266 5296
rect 189718 5176 189724 5228
rect 189776 5216 189782 5228
rect 282914 5216 282920 5228
rect 189776 5188 282920 5216
rect 189776 5176 189782 5188
rect 282914 5176 282920 5188
rect 282972 5176 282978 5228
rect 327994 5176 328000 5228
rect 328052 5216 328058 5228
rect 367002 5216 367008 5228
rect 328052 5188 367008 5216
rect 328052 5176 328058 5188
rect 367002 5176 367008 5188
rect 367060 5176 367066 5228
rect 372522 5176 372528 5228
rect 372580 5216 372586 5228
rect 540790 5216 540796 5228
rect 372580 5188 540796 5216
rect 372580 5176 372586 5188
rect 540790 5176 540796 5188
rect 540848 5176 540854 5228
rect 186130 5108 186136 5160
rect 186188 5148 186194 5160
rect 281534 5148 281540 5160
rect 186188 5120 281540 5148
rect 186188 5108 186194 5120
rect 281534 5108 281540 5120
rect 281592 5108 281598 5160
rect 328178 5108 328184 5160
rect 328236 5148 328242 5160
rect 368198 5148 368204 5160
rect 328236 5120 368204 5148
rect 328236 5108 328242 5120
rect 368198 5108 368204 5120
rect 368256 5108 368262 5160
rect 373902 5108 373908 5160
rect 373960 5148 373966 5160
rect 544378 5148 544384 5160
rect 373960 5120 544384 5148
rect 373960 5108 373966 5120
rect 544378 5108 544384 5120
rect 544436 5108 544442 5160
rect 182542 5040 182548 5092
rect 182600 5080 182606 5092
rect 280246 5080 280252 5092
rect 182600 5052 280252 5080
rect 182600 5040 182606 5052
rect 280246 5040 280252 5052
rect 280304 5040 280310 5092
rect 329650 5040 329656 5092
rect 329708 5080 329714 5092
rect 370590 5080 370596 5092
rect 329708 5052 370596 5080
rect 329708 5040 329714 5052
rect 370590 5040 370596 5052
rect 370648 5040 370654 5092
rect 373810 5040 373816 5092
rect 373868 5080 373874 5092
rect 547874 5080 547880 5092
rect 373868 5052 547880 5080
rect 373868 5040 373874 5052
rect 547874 5040 547880 5052
rect 547932 5040 547938 5092
rect 179046 4972 179052 5024
rect 179104 5012 179110 5024
rect 280154 5012 280160 5024
rect 179104 4984 280160 5012
rect 179104 4972 179110 4984
rect 280154 4972 280160 4984
rect 280212 4972 280218 5024
rect 329466 4972 329472 5024
rect 329524 5012 329530 5024
rect 371694 5012 371700 5024
rect 329524 4984 371700 5012
rect 329524 4972 329530 4984
rect 371694 4972 371700 4984
rect 371752 4972 371758 5024
rect 375006 4972 375012 5024
rect 375064 5012 375070 5024
rect 551462 5012 551468 5024
rect 375064 4984 551468 5012
rect 375064 4972 375070 4984
rect 551462 4972 551468 4984
rect 551520 4972 551526 5024
rect 7650 4904 7656 4956
rect 7708 4944 7714 4956
rect 234525 4947 234583 4953
rect 234525 4944 234537 4947
rect 7708 4916 234537 4944
rect 7708 4904 7714 4916
rect 234525 4913 234537 4916
rect 234571 4913 234583 4947
rect 234525 4907 234583 4913
rect 234614 4904 234620 4956
rect 234672 4944 234678 4956
rect 244829 4947 244887 4953
rect 244829 4944 244841 4947
rect 234672 4916 244841 4944
rect 234672 4904 234678 4916
rect 244829 4913 244841 4916
rect 244875 4913 244887 4947
rect 244829 4907 244887 4913
rect 244936 4916 248414 4944
rect 2866 4836 2872 4888
rect 2924 4876 2930 4888
rect 234706 4876 234712 4888
rect 2924 4848 234712 4876
rect 2924 4836 2930 4848
rect 234706 4836 234712 4848
rect 234764 4836 234770 4888
rect 234801 4879 234859 4885
rect 234801 4845 234813 4879
rect 234847 4876 234859 4879
rect 236086 4876 236092 4888
rect 234847 4848 236092 4876
rect 234847 4845 234859 4848
rect 234801 4839 234859 4845
rect 236086 4836 236092 4848
rect 236144 4836 236150 4888
rect 237006 4836 237012 4888
rect 237064 4876 237070 4888
rect 244936 4876 244964 4916
rect 237064 4848 244964 4876
rect 248386 4876 248414 4916
rect 271230 4904 271236 4956
rect 271288 4944 271294 4956
rect 302418 4944 302424 4956
rect 271288 4916 302424 4944
rect 271288 4904 271294 4916
rect 302418 4904 302424 4916
rect 302476 4904 302482 4956
rect 329558 4904 329564 4956
rect 329616 4944 329622 4956
rect 374086 4944 374092 4956
rect 329616 4916 374092 4944
rect 329616 4904 329622 4916
rect 374086 4904 374092 4916
rect 374144 4904 374150 4956
rect 375098 4904 375104 4956
rect 375156 4944 375162 4956
rect 554958 4944 554964 4956
rect 375156 4916 554964 4944
rect 375156 4904 375162 4916
rect 554958 4904 554964 4916
rect 555016 4904 555022 4956
rect 294046 4876 294052 4888
rect 248386 4848 294052 4876
rect 237064 4836 237070 4848
rect 294046 4836 294052 4848
rect 294104 4836 294110 4888
rect 330846 4836 330852 4888
rect 330904 4876 330910 4888
rect 377674 4876 377680 4888
rect 330904 4848 377680 4876
rect 330904 4836 330910 4848
rect 377674 4836 377680 4848
rect 377732 4836 377738 4888
rect 378042 4836 378048 4888
rect 378100 4876 378106 4888
rect 562042 4876 562048 4888
rect 378100 4848 562048 4876
rect 378100 4836 378106 4848
rect 562042 4836 562048 4848
rect 562100 4836 562106 4888
rect 1670 4768 1676 4820
rect 1728 4808 1734 4820
rect 231949 4811 232007 4817
rect 231949 4808 231961 4811
rect 1728 4780 231961 4808
rect 1728 4768 1734 4780
rect 231949 4777 231961 4780
rect 231995 4777 232007 4811
rect 231949 4771 232007 4777
rect 232222 4768 232228 4820
rect 232280 4808 232286 4820
rect 243541 4811 243599 4817
rect 243541 4808 243553 4811
rect 232280 4780 243553 4808
rect 232280 4768 232286 4780
rect 243541 4777 243553 4780
rect 243587 4777 243599 4811
rect 243541 4771 243599 4777
rect 243633 4811 243691 4817
rect 243633 4777 243645 4811
rect 243679 4808 243691 4811
rect 244918 4808 244924 4820
rect 243679 4780 244924 4808
rect 243679 4777 243691 4780
rect 243633 4771 243691 4777
rect 244918 4768 244924 4780
rect 244976 4768 244982 4820
rect 245013 4811 245071 4817
rect 245013 4777 245025 4811
rect 245059 4808 245071 4811
rect 294138 4808 294144 4820
rect 245059 4780 294144 4808
rect 245059 4777 245071 4780
rect 245013 4771 245071 4777
rect 294138 4768 294144 4780
rect 294196 4768 294202 4820
rect 330754 4768 330760 4820
rect 330812 4808 330818 4820
rect 378870 4808 378876 4820
rect 330812 4780 378876 4808
rect 330812 4768 330818 4780
rect 378870 4768 378876 4780
rect 378928 4768 378934 4820
rect 379330 4768 379336 4820
rect 379388 4808 379394 4820
rect 569126 4808 569132 4820
rect 379388 4780 569132 4808
rect 379388 4768 379394 4780
rect 569126 4768 569132 4780
rect 569184 4768 569190 4820
rect 207382 4700 207388 4752
rect 207440 4740 207446 4752
rect 287054 4740 287060 4752
rect 207440 4712 287060 4740
rect 207440 4700 207446 4712
rect 287054 4700 287060 4712
rect 287112 4700 287118 4752
rect 325418 4700 325424 4752
rect 325476 4740 325482 4752
rect 357526 4740 357532 4752
rect 325476 4712 357532 4740
rect 325476 4700 325482 4712
rect 357526 4700 357532 4712
rect 357584 4700 357590 4752
rect 368290 4700 368296 4752
rect 368348 4740 368354 4752
rect 523034 4740 523040 4752
rect 368348 4712 523040 4740
rect 368348 4700 368354 4712
rect 523034 4700 523040 4712
rect 523092 4700 523098 4752
rect 210970 4632 210976 4684
rect 211028 4672 211034 4684
rect 287146 4672 287152 4684
rect 211028 4644 287152 4672
rect 211028 4632 211034 4644
rect 287146 4632 287152 4644
rect 287204 4632 287210 4684
rect 325510 4632 325516 4684
rect 325568 4672 325574 4684
rect 356330 4672 356336 4684
rect 325568 4644 356336 4672
rect 325568 4632 325574 4644
rect 356330 4632 356336 4644
rect 356388 4632 356394 4684
rect 366910 4632 366916 4684
rect 366968 4672 366974 4684
rect 519538 4672 519544 4684
rect 366968 4644 519544 4672
rect 366968 4632 366974 4644
rect 519538 4632 519544 4644
rect 519596 4632 519602 4684
rect 214466 4564 214472 4616
rect 214524 4604 214530 4616
rect 288434 4604 288440 4616
rect 214524 4576 288440 4604
rect 214524 4564 214530 4576
rect 288434 4564 288440 4576
rect 288492 4564 288498 4616
rect 325326 4564 325332 4616
rect 325384 4604 325390 4616
rect 354030 4604 354036 4616
rect 325384 4576 354036 4604
rect 325384 4564 325390 4576
rect 354030 4564 354036 4576
rect 354088 4564 354094 4616
rect 365622 4564 365628 4616
rect 365680 4604 365686 4616
rect 515950 4604 515956 4616
rect 365680 4576 515956 4604
rect 365680 4564 365686 4576
rect 515950 4564 515956 4576
rect 516008 4564 516014 4616
rect 171962 4496 171968 4548
rect 172020 4536 172026 4548
rect 245010 4536 245016 4548
rect 172020 4508 245016 4536
rect 172020 4496 172026 4508
rect 245010 4496 245016 4508
rect 245068 4496 245074 4548
rect 274818 4496 274824 4548
rect 274876 4536 274882 4548
rect 303798 4536 303804 4548
rect 274876 4508 303804 4536
rect 274876 4496 274882 4508
rect 303798 4496 303804 4508
rect 303856 4496 303862 4548
rect 323946 4496 323952 4548
rect 324004 4536 324010 4548
rect 352834 4536 352840 4548
rect 324004 4508 352840 4536
rect 324004 4496 324010 4508
rect 352834 4496 352840 4508
rect 352892 4496 352898 4548
rect 365530 4496 365536 4548
rect 365588 4536 365594 4548
rect 512454 4536 512460 4548
rect 365588 4508 512460 4536
rect 365588 4496 365594 4508
rect 512454 4496 512460 4508
rect 512512 4496 512518 4548
rect 221550 4428 221556 4480
rect 221608 4468 221614 4480
rect 290090 4468 290096 4480
rect 221608 4440 290096 4468
rect 221608 4428 221614 4440
rect 290090 4428 290096 4440
rect 290148 4428 290154 4480
rect 323854 4428 323860 4480
rect 323912 4468 323918 4480
rect 349246 4468 349252 4480
rect 323912 4440 349252 4468
rect 323912 4428 323918 4440
rect 349246 4428 349252 4440
rect 349304 4428 349310 4480
rect 364242 4428 364248 4480
rect 364300 4468 364306 4480
rect 508866 4468 508872 4480
rect 364300 4440 508872 4468
rect 364300 4428 364306 4440
rect 508866 4428 508872 4440
rect 508924 4428 508930 4480
rect 225138 4360 225144 4412
rect 225196 4400 225202 4412
rect 291194 4400 291200 4412
rect 225196 4372 291200 4400
rect 225196 4360 225202 4372
rect 291194 4360 291200 4372
rect 291252 4360 291258 4412
rect 322658 4360 322664 4412
rect 322716 4400 322722 4412
rect 345750 4400 345756 4412
rect 322716 4372 345756 4400
rect 322716 4360 322722 4372
rect 345750 4360 345756 4372
rect 345808 4360 345814 4412
rect 362770 4360 362776 4412
rect 362828 4400 362834 4412
rect 505370 4400 505376 4412
rect 362828 4372 505376 4400
rect 362828 4360 362834 4372
rect 505370 4360 505376 4372
rect 505428 4360 505434 4412
rect 228726 4292 228732 4344
rect 228784 4332 228790 4344
rect 292666 4332 292672 4344
rect 228784 4304 292672 4332
rect 228784 4292 228790 4304
rect 292666 4292 292672 4304
rect 292724 4292 292730 4344
rect 362862 4292 362868 4344
rect 362920 4332 362926 4344
rect 501782 4332 501788 4344
rect 362920 4304 501788 4332
rect 362920 4292 362926 4304
rect 501782 4292 501788 4304
rect 501840 4292 501846 4344
rect 231949 4267 232007 4273
rect 231949 4233 231961 4267
rect 231995 4264 232007 4267
rect 234798 4264 234804 4276
rect 231995 4236 234804 4264
rect 231995 4233 232007 4236
rect 231949 4227 232007 4233
rect 234798 4224 234804 4236
rect 234856 4224 234862 4276
rect 235810 4224 235816 4276
rect 235868 4264 235874 4276
rect 240137 4267 240195 4273
rect 240137 4264 240149 4267
rect 235868 4236 240149 4264
rect 235868 4224 235874 4236
rect 240137 4233 240149 4236
rect 240183 4233 240195 4267
rect 243449 4267 243507 4273
rect 243449 4264 243461 4267
rect 240137 4227 240195 4233
rect 240244 4236 243461 4264
rect 143534 4156 143540 4208
rect 143592 4196 143598 4208
rect 144822 4196 144828 4208
rect 143592 4168 144828 4196
rect 143592 4156 143598 4168
rect 144822 4156 144828 4168
rect 144880 4156 144886 4208
rect 218054 4156 218060 4208
rect 218112 4196 218118 4208
rect 240244 4196 240272 4236
rect 243449 4233 243461 4236
rect 243495 4233 243507 4267
rect 243449 4227 243507 4233
rect 243541 4267 243599 4273
rect 243541 4233 243553 4267
rect 243587 4264 243599 4267
rect 292574 4264 292580 4276
rect 243587 4236 292580 4264
rect 243587 4233 243599 4236
rect 243541 4227 243599 4233
rect 292574 4224 292580 4236
rect 292632 4224 292638 4276
rect 361482 4224 361488 4276
rect 361540 4264 361546 4276
rect 498194 4264 498200 4276
rect 361540 4236 498200 4264
rect 361540 4224 361546 4236
rect 498194 4224 498200 4236
rect 498252 4224 498258 4276
rect 218112 4168 240272 4196
rect 240321 4199 240379 4205
rect 218112 4156 218118 4168
rect 240321 4165 240333 4199
rect 240367 4196 240379 4199
rect 293954 4196 293960 4208
rect 240367 4168 293960 4196
rect 240367 4165 240379 4168
rect 240321 4159 240379 4165
rect 293954 4156 293960 4168
rect 294012 4156 294018 4208
rect 332410 4156 332416 4208
rect 332468 4196 332474 4208
rect 381170 4196 381176 4208
rect 332468 4168 381176 4196
rect 332468 4156 332474 4168
rect 381170 4156 381176 4168
rect 381228 4156 381234 4208
rect 489914 4156 489920 4208
rect 489972 4196 489978 4208
rect 491110 4196 491116 4208
rect 489972 4168 491116 4196
rect 489972 4156 489978 4168
rect 491110 4156 491116 4168
rect 491168 4156 491174 4208
rect 50154 4088 50160 4140
rect 50212 4128 50218 4140
rect 241517 4131 241575 4137
rect 241517 4128 241529 4131
rect 50212 4100 241529 4128
rect 50212 4088 50218 4100
rect 241517 4097 241529 4100
rect 241563 4097 241575 4131
rect 245930 4128 245936 4140
rect 241517 4091 241575 4097
rect 241624 4100 245936 4128
rect 46658 4020 46664 4072
rect 46716 4060 46722 4072
rect 241624 4060 241652 4100
rect 245930 4088 245936 4100
rect 245988 4088 245994 4140
rect 279510 4088 279516 4140
rect 279568 4128 279574 4140
rect 305270 4128 305276 4140
rect 279568 4100 305276 4128
rect 279568 4088 279574 4100
rect 305270 4088 305276 4100
rect 305328 4088 305334 4140
rect 305365 4131 305423 4137
rect 305365 4097 305377 4131
rect 305411 4128 305423 4131
rect 307938 4128 307944 4140
rect 305411 4100 307944 4128
rect 305411 4097 305423 4100
rect 305365 4091 305423 4097
rect 307938 4088 307944 4100
rect 307996 4088 308002 4140
rect 328362 4088 328368 4140
rect 328420 4128 328426 4140
rect 331677 4131 331735 4137
rect 331677 4128 331689 4131
rect 328420 4100 331689 4128
rect 328420 4088 328426 4100
rect 331677 4097 331689 4100
rect 331723 4097 331735 4131
rect 331677 4091 331735 4097
rect 332502 4088 332508 4140
rect 332560 4128 332566 4140
rect 334069 4131 334127 4137
rect 332560 4100 334020 4128
rect 332560 4088 332566 4100
rect 46716 4032 241652 4060
rect 46716 4020 46722 4032
rect 244090 4020 244096 4072
rect 244148 4060 244154 4072
rect 249058 4060 249064 4072
rect 244148 4032 249064 4060
rect 244148 4020 244154 4032
rect 249058 4020 249064 4032
rect 249116 4020 249122 4072
rect 276014 4020 276020 4072
rect 276072 4060 276078 4072
rect 303890 4060 303896 4072
rect 276072 4032 303896 4060
rect 276072 4020 276078 4032
rect 303890 4020 303896 4032
rect 303948 4020 303954 4072
rect 320082 4020 320088 4072
rect 320140 4060 320146 4072
rect 333882 4060 333888 4072
rect 320140 4032 333888 4060
rect 320140 4020 320146 4032
rect 333882 4020 333888 4032
rect 333940 4020 333946 4072
rect 333992 4069 334020 4100
rect 334069 4097 334081 4131
rect 334115 4128 334127 4131
rect 365806 4128 365812 4140
rect 334115 4100 365812 4128
rect 334115 4097 334127 4100
rect 334069 4091 334127 4097
rect 365806 4088 365812 4100
rect 365864 4088 365870 4140
rect 396718 4088 396724 4140
rect 396776 4128 396782 4140
rect 521838 4128 521844 4140
rect 396776 4100 521844 4128
rect 396776 4088 396782 4100
rect 521838 4088 521844 4100
rect 521896 4088 521902 4140
rect 333977 4063 334035 4069
rect 333977 4029 333989 4063
rect 334023 4029 334035 4063
rect 376478 4060 376484 4072
rect 333977 4023 334035 4029
rect 334084 4032 376484 4060
rect 45370 3952 45376 4004
rect 45428 3992 45434 4004
rect 245746 3992 245752 4004
rect 45428 3964 245752 3992
rect 45428 3952 45434 3964
rect 245746 3952 245752 3964
rect 245804 3952 245810 4004
rect 277118 3952 277124 4004
rect 277176 3992 277182 4004
rect 305086 3992 305092 4004
rect 277176 3964 305092 3992
rect 277176 3952 277182 3964
rect 305086 3952 305092 3964
rect 305144 3952 305150 4004
rect 324958 3952 324964 4004
rect 325016 3992 325022 4004
rect 332686 3992 332692 4004
rect 325016 3964 332692 3992
rect 325016 3952 325022 3964
rect 332686 3952 332692 3964
rect 332744 3952 332750 4004
rect 39574 3884 39580 3936
rect 39632 3924 39638 3936
rect 244366 3924 244372 3936
rect 39632 3896 244372 3924
rect 39632 3884 39638 3896
rect 244366 3884 244372 3896
rect 244424 3884 244430 3936
rect 265342 3884 265348 3936
rect 265400 3924 265406 3936
rect 271138 3924 271144 3936
rect 265400 3896 271144 3924
rect 265400 3884 265406 3896
rect 271138 3884 271144 3896
rect 271196 3884 271202 3936
rect 272426 3884 272432 3936
rect 272484 3924 272490 3936
rect 303706 3924 303712 3936
rect 272484 3896 303712 3924
rect 272484 3884 272490 3896
rect 303706 3884 303712 3896
rect 303764 3884 303770 3936
rect 305546 3884 305552 3936
rect 305604 3924 305610 3936
rect 311986 3924 311992 3936
rect 305604 3896 311992 3924
rect 305604 3884 305610 3896
rect 311986 3884 311992 3896
rect 312044 3884 312050 3936
rect 326982 3884 326988 3936
rect 327040 3924 327046 3936
rect 330573 3927 330631 3933
rect 330573 3924 330585 3927
rect 327040 3896 330585 3924
rect 327040 3884 327046 3896
rect 330573 3893 330585 3896
rect 330619 3893 330631 3927
rect 330573 3887 330631 3893
rect 331122 3884 331128 3936
rect 331180 3924 331186 3936
rect 334084 3924 334112 4032
rect 376478 4020 376484 4032
rect 376536 4020 376542 4072
rect 399478 4020 399484 4072
rect 399536 4060 399542 4072
rect 529014 4060 529020 4072
rect 399536 4032 529020 4060
rect 399536 4020 399542 4032
rect 529014 4020 529020 4032
rect 529072 4020 529078 4072
rect 334253 3995 334311 4001
rect 334253 3961 334265 3995
rect 334299 3992 334311 3995
rect 336921 3995 336979 4001
rect 334299 3964 336872 3992
rect 334299 3961 334311 3964
rect 334253 3955 334311 3961
rect 331180 3896 334112 3924
rect 334161 3927 334219 3933
rect 331180 3884 331186 3896
rect 334161 3893 334173 3927
rect 334207 3924 334219 3927
rect 336737 3927 336795 3933
rect 336737 3924 336749 3927
rect 334207 3896 336749 3924
rect 334207 3893 334219 3896
rect 334161 3887 334219 3893
rect 336737 3893 336749 3896
rect 336783 3893 336795 3927
rect 336844 3924 336872 3964
rect 336921 3961 336933 3995
rect 336967 3992 336979 3995
rect 379974 3992 379980 4004
rect 336967 3964 379980 3992
rect 336967 3961 336979 3964
rect 336921 3955 336979 3961
rect 379974 3952 379980 3964
rect 380032 3952 380038 4004
rect 404998 3952 405004 4004
rect 405056 3992 405062 4004
rect 536098 3992 536104 4004
rect 405056 3964 536104 3992
rect 405056 3952 405062 3964
rect 536098 3952 536104 3964
rect 536156 3952 536162 4004
rect 383562 3924 383568 3936
rect 336844 3896 383568 3924
rect 336737 3887 336795 3893
rect 383562 3884 383568 3896
rect 383620 3884 383626 3936
rect 403618 3884 403624 3936
rect 403676 3924 403682 3936
rect 543182 3924 543188 3936
rect 403676 3896 543188 3924
rect 403676 3884 403682 3896
rect 543182 3884 543188 3896
rect 543240 3884 543246 3936
rect 35986 3816 35992 3868
rect 36044 3856 36050 3868
rect 37090 3856 37096 3868
rect 36044 3828 37096 3856
rect 36044 3816 36050 3828
rect 37090 3816 37096 3828
rect 37148 3816 37154 3868
rect 38378 3816 38384 3868
rect 38436 3856 38442 3868
rect 244642 3856 244648 3868
rect 38436 3828 244648 3856
rect 38436 3816 38442 3828
rect 244642 3816 244648 3828
rect 244700 3816 244706 3868
rect 270034 3816 270040 3868
rect 270092 3856 270098 3868
rect 302326 3856 302332 3868
rect 270092 3828 302332 3856
rect 270092 3816 270098 3828
rect 302326 3816 302332 3828
rect 302384 3816 302390 3868
rect 304350 3816 304356 3868
rect 304408 3856 304414 3868
rect 311158 3856 311164 3868
rect 304408 3828 311164 3856
rect 304408 3816 304414 3828
rect 311158 3816 311164 3828
rect 311216 3816 311222 3868
rect 320818 3816 320824 3868
rect 320876 3856 320882 3868
rect 326798 3856 326804 3868
rect 320876 3828 326804 3856
rect 320876 3816 320882 3828
rect 326798 3816 326804 3828
rect 326856 3816 326862 3868
rect 328270 3816 328276 3868
rect 328328 3856 328334 3868
rect 333701 3859 333759 3865
rect 333701 3856 333713 3859
rect 328328 3828 333713 3856
rect 328328 3816 328334 3828
rect 333701 3825 333713 3828
rect 333747 3825 333759 3859
rect 333701 3819 333759 3825
rect 333790 3816 333796 3868
rect 333848 3856 333854 3868
rect 387150 3856 387156 3868
rect 333848 3828 387156 3856
rect 333848 3816 333854 3828
rect 387150 3816 387156 3828
rect 387208 3816 387214 3868
rect 411898 3816 411904 3868
rect 411956 3856 411962 3868
rect 557350 3856 557356 3868
rect 411956 3828 557356 3856
rect 411956 3816 411962 3828
rect 557350 3816 557356 3828
rect 557408 3816 557414 3868
rect 31294 3748 31300 3800
rect 31352 3788 31358 3800
rect 241882 3788 241888 3800
rect 31352 3760 241888 3788
rect 31352 3748 31358 3760
rect 241882 3748 241888 3760
rect 241940 3748 241946 3800
rect 264146 3748 264152 3800
rect 264204 3788 264210 3800
rect 301130 3788 301136 3800
rect 264204 3760 301136 3788
rect 264204 3748 264210 3760
rect 301130 3748 301136 3760
rect 301188 3748 301194 3800
rect 301958 3748 301964 3800
rect 302016 3788 302022 3800
rect 310790 3788 310796 3800
rect 302016 3760 310796 3788
rect 302016 3748 302022 3760
rect 310790 3748 310796 3760
rect 310848 3748 310854 3800
rect 322198 3748 322204 3800
rect 322256 3788 322262 3800
rect 330386 3788 330392 3800
rect 322256 3760 330392 3788
rect 322256 3748 322262 3760
rect 330386 3748 330392 3760
rect 330444 3748 330450 3800
rect 342162 3788 342168 3800
rect 330496 3760 342168 3788
rect 32398 3680 32404 3732
rect 32456 3720 32462 3732
rect 243078 3720 243084 3732
rect 32456 3692 243084 3720
rect 32456 3680 32462 3692
rect 243078 3680 243084 3692
rect 243136 3680 243142 3732
rect 245194 3680 245200 3732
rect 245252 3720 245258 3732
rect 254578 3720 254584 3732
rect 245252 3692 254584 3720
rect 245252 3680 245258 3692
rect 254578 3680 254584 3692
rect 254636 3680 254642 3732
rect 257062 3680 257068 3732
rect 257120 3720 257126 3732
rect 299658 3720 299664 3732
rect 257120 3692 299664 3720
rect 257120 3680 257126 3692
rect 299658 3680 299664 3692
rect 299716 3680 299722 3732
rect 301041 3723 301099 3729
rect 301041 3689 301053 3723
rect 301087 3720 301099 3723
rect 305454 3720 305460 3732
rect 301087 3692 305460 3720
rect 301087 3689 301099 3692
rect 301041 3683 301099 3689
rect 305454 3680 305460 3692
rect 305512 3680 305518 3732
rect 306469 3723 306527 3729
rect 306469 3689 306481 3723
rect 306515 3720 306527 3723
rect 310698 3720 310704 3732
rect 306515 3692 310704 3720
rect 306515 3689 306527 3692
rect 306469 3683 306527 3689
rect 310698 3680 310704 3692
rect 310756 3680 310762 3732
rect 321278 3680 321284 3732
rect 321336 3720 321342 3732
rect 330496 3720 330524 3760
rect 342162 3748 342168 3760
rect 342220 3748 342226 3800
rect 343542 3748 343548 3800
rect 343600 3788 343606 3800
rect 426158 3788 426164 3800
rect 343600 3760 426164 3788
rect 343600 3748 343606 3760
rect 426158 3748 426164 3760
rect 426216 3748 426222 3800
rect 429749 3791 429807 3797
rect 429749 3788 429761 3791
rect 426268 3760 429761 3788
rect 321336 3692 330524 3720
rect 330573 3723 330631 3729
rect 321336 3680 321342 3692
rect 330573 3689 330585 3723
rect 330619 3720 330631 3723
rect 333609 3723 333667 3729
rect 333609 3720 333621 3723
rect 330619 3692 333621 3720
rect 330619 3689 330631 3692
rect 330573 3683 330631 3689
rect 333609 3689 333621 3692
rect 333655 3689 333667 3723
rect 333609 3683 333667 3689
rect 333698 3680 333704 3732
rect 333756 3720 333762 3732
rect 390646 3720 390652 3732
rect 333756 3692 390652 3720
rect 333756 3680 333762 3692
rect 390646 3680 390652 3692
rect 390704 3680 390710 3732
rect 391198 3680 391204 3732
rect 391256 3720 391262 3732
rect 415486 3720 415492 3732
rect 391256 3692 415492 3720
rect 391256 3680 391262 3692
rect 415486 3680 415492 3692
rect 415544 3680 415550 3732
rect 416038 3680 416044 3732
rect 416096 3720 416102 3732
rect 422570 3720 422576 3732
rect 416096 3692 422576 3720
rect 416096 3680 416102 3692
rect 422570 3680 422576 3692
rect 422628 3680 422634 3732
rect 425698 3680 425704 3732
rect 425756 3720 425762 3732
rect 426268 3720 426296 3760
rect 429749 3757 429761 3760
rect 429795 3757 429807 3791
rect 429749 3751 429807 3757
rect 429838 3748 429844 3800
rect 429896 3788 429902 3800
rect 432506 3788 432512 3800
rect 429896 3760 432512 3788
rect 429896 3748 429902 3760
rect 432506 3748 432512 3760
rect 432564 3748 432570 3800
rect 432598 3748 432604 3800
rect 432656 3788 432662 3800
rect 440326 3788 440332 3800
rect 432656 3760 440332 3788
rect 432656 3748 432662 3760
rect 440326 3748 440332 3760
rect 440384 3748 440390 3800
rect 440421 3791 440479 3797
rect 440421 3757 440433 3791
rect 440467 3788 440479 3791
rect 571518 3788 571524 3800
rect 440467 3760 571524 3788
rect 440467 3757 440479 3760
rect 440421 3751 440479 3757
rect 571518 3748 571524 3760
rect 571576 3748 571582 3800
rect 425756 3692 426296 3720
rect 427081 3723 427139 3729
rect 425756 3680 425762 3692
rect 427081 3689 427093 3723
rect 427127 3720 427139 3723
rect 564434 3720 564440 3732
rect 427127 3692 564440 3720
rect 427127 3689 427139 3692
rect 427081 3683 427139 3689
rect 564434 3680 564440 3692
rect 564492 3680 564498 3732
rect 28810 3612 28816 3664
rect 28868 3652 28874 3664
rect 241606 3652 241612 3664
rect 28868 3624 241612 3652
rect 28868 3612 28874 3624
rect 241606 3612 241612 3624
rect 241664 3612 241670 3664
rect 241698 3612 241704 3664
rect 241756 3652 241762 3664
rect 251818 3652 251824 3664
rect 241756 3624 251824 3652
rect 241756 3612 241762 3624
rect 251818 3612 251824 3624
rect 251876 3612 251882 3664
rect 253474 3612 253480 3664
rect 253532 3652 253538 3664
rect 298462 3652 298468 3664
rect 253532 3624 298468 3652
rect 253532 3612 253538 3624
rect 298462 3612 298468 3624
rect 298520 3612 298526 3664
rect 298554 3612 298560 3664
rect 298612 3652 298618 3664
rect 309134 3652 309140 3664
rect 298612 3624 309140 3652
rect 298612 3612 298618 3624
rect 309134 3612 309140 3624
rect 309192 3612 309198 3664
rect 321370 3612 321376 3664
rect 321428 3652 321434 3664
rect 337470 3652 337476 3664
rect 321428 3624 337476 3652
rect 321428 3612 321434 3624
rect 337470 3612 337476 3624
rect 337528 3612 337534 3664
rect 338758 3612 338764 3664
rect 338816 3652 338822 3664
rect 404814 3652 404820 3664
rect 338816 3624 404820 3652
rect 338816 3612 338822 3624
rect 404814 3612 404820 3624
rect 404872 3612 404878 3664
rect 413278 3612 413284 3664
rect 413336 3652 413342 3664
rect 560846 3652 560852 3664
rect 413336 3624 560852 3652
rect 413336 3612 413342 3624
rect 560846 3612 560852 3624
rect 560904 3612 560910 3664
rect 11146 3544 11152 3596
rect 11204 3584 11210 3596
rect 12342 3584 12348 3596
rect 11204 3556 12348 3584
rect 11204 3544 11210 3556
rect 12342 3544 12348 3556
rect 12400 3544 12406 3596
rect 25314 3544 25320 3596
rect 25372 3584 25378 3596
rect 240502 3584 240508 3596
rect 25372 3556 240508 3584
rect 25372 3544 25378 3556
rect 240502 3544 240508 3556
rect 240560 3544 240566 3596
rect 241517 3587 241575 3593
rect 241517 3553 241529 3587
rect 241563 3584 241575 3587
rect 247034 3584 247040 3596
rect 241563 3556 247040 3584
rect 241563 3553 241575 3556
rect 241517 3547 241575 3553
rect 247034 3544 247040 3556
rect 247092 3544 247098 3596
rect 255866 3544 255872 3596
rect 255924 3584 255930 3596
rect 256602 3584 256608 3596
rect 255924 3556 256608 3584
rect 255924 3544 255930 3556
rect 256602 3544 256608 3556
rect 256660 3544 256666 3596
rect 256697 3587 256755 3593
rect 256697 3553 256709 3587
rect 256743 3584 256755 3587
rect 298186 3584 298192 3596
rect 256743 3556 298192 3584
rect 256743 3553 256755 3556
rect 256697 3547 256755 3553
rect 298186 3544 298192 3556
rect 298244 3544 298250 3596
rect 300762 3544 300768 3596
rect 300820 3584 300826 3596
rect 306469 3587 306527 3593
rect 306469 3584 306481 3587
rect 300820 3556 306481 3584
rect 300820 3544 300826 3556
rect 306469 3553 306481 3556
rect 306515 3553 306527 3587
rect 309318 3584 309324 3596
rect 306469 3547 306527 3553
rect 306576 3556 309324 3584
rect 566 3476 572 3528
rect 624 3516 630 3528
rect 1302 3516 1308 3528
rect 624 3488 1308 3516
rect 624 3476 630 3488
rect 1302 3476 1308 3488
rect 1360 3476 1366 3528
rect 9950 3476 9956 3528
rect 10008 3516 10014 3528
rect 10962 3516 10968 3528
rect 10008 3488 10968 3516
rect 10008 3476 10014 3488
rect 10962 3476 10968 3488
rect 11020 3476 11026 3528
rect 18230 3476 18236 3528
rect 18288 3516 18294 3528
rect 19242 3516 19248 3528
rect 18288 3488 19248 3516
rect 18288 3476 18294 3488
rect 19242 3476 19248 3488
rect 19300 3476 19306 3528
rect 24210 3476 24216 3528
rect 24268 3516 24274 3528
rect 240318 3516 240324 3528
rect 24268 3488 240324 3516
rect 24268 3476 24274 3488
rect 240318 3476 240324 3488
rect 240376 3476 240382 3528
rect 246390 3476 246396 3528
rect 246448 3516 246454 3528
rect 296990 3516 296996 3528
rect 246448 3488 296996 3516
rect 246448 3476 246454 3488
rect 296990 3476 296996 3488
rect 297048 3476 297054 3528
rect 297266 3476 297272 3528
rect 297324 3516 297330 3528
rect 306576 3516 306604 3556
rect 309318 3544 309324 3556
rect 309376 3544 309382 3596
rect 317322 3544 317328 3596
rect 317380 3584 317386 3596
rect 325510 3584 325516 3596
rect 317380 3556 325516 3584
rect 317380 3544 317386 3556
rect 325510 3544 325516 3556
rect 325568 3544 325574 3596
rect 327718 3544 327724 3596
rect 327776 3584 327782 3596
rect 331582 3584 331588 3596
rect 327776 3556 331588 3584
rect 327776 3544 327782 3556
rect 331582 3544 331588 3556
rect 331640 3544 331646 3596
rect 331677 3587 331735 3593
rect 331677 3553 331689 3587
rect 331723 3584 331735 3587
rect 369394 3584 369400 3596
rect 331723 3556 369400 3584
rect 331723 3553 331735 3556
rect 331677 3547 331735 3553
rect 369394 3544 369400 3556
rect 369452 3544 369458 3596
rect 369762 3544 369768 3596
rect 369820 3584 369826 3596
rect 532510 3584 532516 3596
rect 369820 3556 532516 3584
rect 369820 3544 369826 3556
rect 532510 3544 532516 3556
rect 532568 3544 532574 3596
rect 297324 3488 306604 3516
rect 297324 3476 297330 3488
rect 306742 3476 306748 3528
rect 306800 3516 306806 3528
rect 307662 3516 307668 3528
rect 306800 3488 307668 3516
rect 306800 3476 306806 3488
rect 307662 3476 307668 3488
rect 307720 3476 307726 3528
rect 309226 3516 309232 3528
rect 307772 3488 309232 3516
rect 23014 3408 23020 3460
rect 23072 3448 23078 3460
rect 240226 3448 240232 3460
rect 23072 3420 240232 3448
rect 23072 3408 23078 3420
rect 240226 3408 240232 3420
rect 240284 3408 240290 3460
rect 242894 3408 242900 3460
rect 242952 3448 242958 3460
rect 242952 3420 277394 3448
rect 242952 3408 242958 3420
rect 27706 3340 27712 3392
rect 27764 3380 27770 3392
rect 28902 3380 28908 3392
rect 27764 3352 28908 3380
rect 27764 3340 27770 3352
rect 28902 3340 28908 3352
rect 28960 3340 28966 3392
rect 34790 3340 34796 3392
rect 34848 3380 34854 3392
rect 35802 3380 35808 3392
rect 34848 3352 35808 3380
rect 34848 3340 34854 3352
rect 35802 3340 35808 3352
rect 35860 3340 35866 3392
rect 40678 3340 40684 3392
rect 40736 3380 40742 3392
rect 41322 3380 41328 3392
rect 40736 3352 41328 3380
rect 40736 3340 40742 3352
rect 41322 3340 41328 3352
rect 41380 3340 41386 3392
rect 41874 3340 41880 3392
rect 41932 3380 41938 3392
rect 42702 3380 42708 3392
rect 41932 3352 42708 3380
rect 41932 3340 41938 3352
rect 42702 3340 42708 3352
rect 42760 3340 42766 3392
rect 43070 3340 43076 3392
rect 43128 3380 43134 3392
rect 44082 3380 44088 3392
rect 43128 3352 44088 3380
rect 43128 3340 43134 3352
rect 44082 3340 44088 3352
rect 44140 3340 44146 3392
rect 44266 3340 44272 3392
rect 44324 3380 44330 3392
rect 45462 3380 45468 3392
rect 44324 3352 45468 3380
rect 44324 3340 44330 3352
rect 45462 3340 45468 3352
rect 45520 3340 45526 3392
rect 48958 3340 48964 3392
rect 49016 3380 49022 3392
rect 49602 3380 49608 3392
rect 49016 3352 49608 3380
rect 49016 3340 49022 3352
rect 49602 3340 49608 3352
rect 49660 3340 49666 3392
rect 52546 3340 52552 3392
rect 52604 3380 52610 3392
rect 53650 3380 53656 3392
rect 52604 3352 53656 3380
rect 52604 3340 52610 3352
rect 53650 3340 53656 3352
rect 53708 3340 53714 3392
rect 56042 3340 56048 3392
rect 56100 3380 56106 3392
rect 56502 3380 56508 3392
rect 56100 3352 56508 3380
rect 56100 3340 56106 3352
rect 56502 3340 56508 3352
rect 56560 3340 56566 3392
rect 59630 3340 59636 3392
rect 59688 3380 59694 3392
rect 60642 3380 60648 3392
rect 59688 3352 60648 3380
rect 59688 3340 59694 3352
rect 60642 3340 60648 3352
rect 60700 3340 60706 3392
rect 60826 3340 60832 3392
rect 60884 3380 60890 3392
rect 62022 3380 62028 3392
rect 60884 3352 62028 3380
rect 60884 3340 60890 3352
rect 62022 3340 62028 3352
rect 62080 3340 62086 3392
rect 66714 3340 66720 3392
rect 66772 3380 66778 3392
rect 67542 3380 67548 3392
rect 66772 3352 67548 3380
rect 66772 3340 66778 3352
rect 67542 3340 67548 3352
rect 67600 3340 67606 3392
rect 67910 3340 67916 3392
rect 67968 3380 67974 3392
rect 68922 3380 68928 3392
rect 67968 3352 68928 3380
rect 67968 3340 67974 3352
rect 68922 3340 68928 3352
rect 68980 3340 68986 3392
rect 248690 3380 248696 3392
rect 69032 3352 248696 3380
rect 57238 3272 57244 3324
rect 57296 3312 57302 3324
rect 69032 3312 69060 3352
rect 248690 3340 248696 3352
rect 248748 3340 248754 3392
rect 249978 3340 249984 3392
rect 250036 3380 250042 3392
rect 256697 3383 256755 3389
rect 256697 3380 256709 3383
rect 250036 3352 256709 3380
rect 250036 3340 250042 3352
rect 256697 3349 256709 3352
rect 256743 3349 256755 3383
rect 256697 3343 256755 3349
rect 259454 3340 259460 3392
rect 259512 3380 259518 3392
rect 260742 3380 260748 3392
rect 259512 3352 260748 3380
rect 259512 3340 259518 3352
rect 260742 3340 260748 3352
rect 260800 3340 260806 3392
rect 273622 3340 273628 3392
rect 273680 3380 273686 3392
rect 274542 3380 274548 3392
rect 273680 3352 274548 3380
rect 273680 3340 273686 3352
rect 274542 3340 274548 3352
rect 274600 3340 274606 3392
rect 277366 3380 277394 3420
rect 278314 3408 278320 3460
rect 278372 3448 278378 3460
rect 282178 3448 282184 3460
rect 278372 3420 282184 3448
rect 278372 3408 278378 3420
rect 282178 3408 282184 3420
rect 282236 3408 282242 3460
rect 284294 3408 284300 3460
rect 284352 3448 284358 3460
rect 285582 3448 285588 3460
rect 284352 3420 285588 3448
rect 284352 3408 284358 3420
rect 285582 3408 285588 3420
rect 285640 3408 285646 3460
rect 287790 3408 287796 3460
rect 287848 3448 287854 3460
rect 288342 3448 288348 3460
rect 287848 3420 288348 3448
rect 287848 3408 287854 3420
rect 288342 3408 288348 3420
rect 288400 3408 288406 3460
rect 288986 3408 288992 3460
rect 289044 3448 289050 3460
rect 289722 3448 289728 3460
rect 289044 3420 289728 3448
rect 289044 3408 289050 3420
rect 289722 3408 289728 3420
rect 289780 3408 289786 3460
rect 295702 3448 295708 3460
rect 289832 3420 295708 3448
rect 289832 3380 289860 3420
rect 295702 3408 295708 3420
rect 295760 3408 295766 3460
rect 296070 3408 296076 3460
rect 296128 3448 296134 3460
rect 307772 3448 307800 3488
rect 309226 3476 309232 3488
rect 309284 3476 309290 3528
rect 313274 3476 313280 3528
rect 313332 3516 313338 3528
rect 313826 3516 313832 3528
rect 313332 3488 313832 3516
rect 313332 3476 313338 3488
rect 313826 3476 313832 3488
rect 313884 3476 313890 3528
rect 320910 3476 320916 3528
rect 320968 3516 320974 3528
rect 322106 3516 322112 3528
rect 320968 3488 322112 3516
rect 320968 3476 320974 3488
rect 322106 3476 322112 3488
rect 322164 3476 322170 3528
rect 322290 3476 322296 3528
rect 322348 3516 322354 3528
rect 323302 3516 323308 3528
rect 322348 3488 323308 3516
rect 322348 3476 322354 3488
rect 323302 3476 323308 3488
rect 323360 3476 323366 3528
rect 327994 3516 328000 3528
rect 323412 3488 328000 3516
rect 296128 3420 307800 3448
rect 296128 3408 296134 3420
rect 309042 3408 309048 3460
rect 309100 3448 309106 3460
rect 312170 3448 312176 3460
rect 309100 3420 312176 3448
rect 309100 3408 309106 3420
rect 312170 3408 312176 3420
rect 312228 3408 312234 3460
rect 277366 3352 289860 3380
rect 290645 3383 290703 3389
rect 290645 3349 290657 3383
rect 290691 3380 290703 3383
rect 299569 3383 299627 3389
rect 299569 3380 299581 3383
rect 290691 3352 299581 3380
rect 290691 3349 290703 3352
rect 290645 3343 290703 3349
rect 299569 3349 299581 3352
rect 299615 3349 299627 3383
rect 299569 3343 299627 3349
rect 299658 3340 299664 3392
rect 299716 3380 299722 3392
rect 299716 3352 306374 3380
rect 299716 3340 299722 3352
rect 251542 3312 251548 3324
rect 57296 3284 69060 3312
rect 69676 3284 251548 3312
rect 57296 3272 57302 3284
rect 64322 3204 64328 3256
rect 64380 3244 64386 3256
rect 69676 3244 69704 3284
rect 251542 3272 251548 3284
rect 251600 3272 251606 3324
rect 283098 3272 283104 3324
rect 283156 3312 283162 3324
rect 301593 3315 301651 3321
rect 283156 3284 301544 3312
rect 283156 3272 283162 3284
rect 64380 3216 69704 3244
rect 64380 3204 64386 3216
rect 73798 3204 73804 3256
rect 73856 3244 73862 3256
rect 74442 3244 74448 3256
rect 73856 3216 74448 3244
rect 73856 3204 73862 3216
rect 74442 3204 74448 3216
rect 74500 3204 74506 3256
rect 74994 3204 75000 3256
rect 75052 3244 75058 3256
rect 75822 3244 75828 3256
rect 75052 3216 75828 3244
rect 75052 3204 75058 3216
rect 75822 3204 75828 3216
rect 75880 3204 75886 3256
rect 77386 3204 77392 3256
rect 77444 3244 77450 3256
rect 78582 3244 78588 3256
rect 77444 3216 78588 3244
rect 77444 3204 77450 3216
rect 78582 3204 78588 3216
rect 78640 3204 78646 3256
rect 80882 3204 80888 3256
rect 80940 3244 80946 3256
rect 81342 3244 81348 3256
rect 80940 3216 81348 3244
rect 80940 3204 80946 3216
rect 81342 3204 81348 3216
rect 81400 3204 81406 3256
rect 82078 3204 82084 3256
rect 82136 3244 82142 3256
rect 82722 3244 82728 3256
rect 82136 3216 82728 3244
rect 82136 3204 82142 3216
rect 82722 3204 82728 3216
rect 82780 3204 82786 3256
rect 84470 3204 84476 3256
rect 84528 3244 84534 3256
rect 85482 3244 85488 3256
rect 84528 3216 85488 3244
rect 84528 3204 84534 3216
rect 85482 3204 85488 3216
rect 85540 3204 85546 3256
rect 85666 3204 85672 3256
rect 85724 3244 85730 3256
rect 86770 3244 86776 3256
rect 85724 3216 86776 3244
rect 85724 3204 85730 3216
rect 86770 3204 86776 3216
rect 86828 3204 86834 3256
rect 90358 3204 90364 3256
rect 90416 3244 90422 3256
rect 91002 3244 91008 3256
rect 90416 3216 91008 3244
rect 90416 3204 90422 3216
rect 91002 3204 91008 3216
rect 91060 3204 91066 3256
rect 91554 3204 91560 3256
rect 91612 3244 91618 3256
rect 92382 3244 92388 3256
rect 91612 3216 92388 3244
rect 91612 3204 91618 3216
rect 92382 3204 92388 3216
rect 92440 3204 92446 3256
rect 252922 3244 252928 3256
rect 92492 3216 252928 3244
rect 71498 3136 71504 3188
rect 71556 3176 71562 3188
rect 92492 3176 92520 3216
rect 252922 3204 252928 3216
rect 252980 3204 252986 3256
rect 281902 3204 281908 3256
rect 281960 3244 281966 3256
rect 301041 3247 301099 3253
rect 301041 3244 301053 3247
rect 281960 3216 301053 3244
rect 281960 3204 281966 3216
rect 301041 3213 301053 3216
rect 301087 3213 301099 3247
rect 301516 3244 301544 3284
rect 301593 3281 301605 3315
rect 301639 3312 301651 3315
rect 305365 3315 305423 3321
rect 305365 3312 305377 3315
rect 301639 3284 305377 3312
rect 301639 3281 301651 3284
rect 301593 3275 301651 3281
rect 305365 3281 305377 3284
rect 305411 3281 305423 3315
rect 306346 3312 306374 3352
rect 307938 3340 307944 3392
rect 307996 3380 308002 3392
rect 312078 3380 312084 3392
rect 307996 3352 312084 3380
rect 307996 3340 308002 3352
rect 312078 3340 312084 3352
rect 312136 3340 312142 3392
rect 318610 3340 318616 3392
rect 318668 3380 318674 3392
rect 323412 3380 323440 3488
rect 327994 3476 328000 3488
rect 328052 3476 328058 3528
rect 331030 3476 331036 3528
rect 331088 3516 331094 3528
rect 334161 3519 334219 3525
rect 334161 3516 334173 3519
rect 331088 3488 334173 3516
rect 331088 3476 331094 3488
rect 334161 3485 334173 3488
rect 334207 3485 334219 3519
rect 334161 3479 334219 3485
rect 334253 3519 334311 3525
rect 334253 3485 334265 3519
rect 334299 3516 334311 3519
rect 372890 3516 372896 3528
rect 334299 3488 372896 3516
rect 334299 3485 334311 3488
rect 334253 3479 334311 3485
rect 372890 3476 372896 3488
rect 372948 3476 372954 3528
rect 375190 3476 375196 3528
rect 375248 3516 375254 3528
rect 550266 3516 550272 3528
rect 375248 3488 550272 3516
rect 375248 3476 375254 3488
rect 550266 3476 550272 3488
rect 550324 3476 550330 3528
rect 324501 3451 324559 3457
rect 324501 3417 324513 3451
rect 324547 3448 324559 3451
rect 329190 3448 329196 3460
rect 324547 3420 329196 3448
rect 324547 3417 324559 3420
rect 324501 3411 324559 3417
rect 329190 3408 329196 3420
rect 329248 3408 329254 3460
rect 330938 3408 330944 3460
rect 330996 3448 331002 3460
rect 375282 3448 375288 3460
rect 330996 3420 375288 3448
rect 330996 3408 331002 3420
rect 375282 3408 375288 3420
rect 375340 3408 375346 3460
rect 375374 3408 375380 3460
rect 375432 3448 375438 3460
rect 553762 3448 553768 3460
rect 375432 3420 553768 3448
rect 375432 3408 375438 3420
rect 553762 3408 553768 3420
rect 553820 3408 553826 3460
rect 318668 3352 323440 3380
rect 318668 3340 318674 3352
rect 324222 3340 324228 3392
rect 324280 3380 324286 3392
rect 351638 3380 351644 3392
rect 324280 3352 351644 3380
rect 324280 3340 324286 3352
rect 351638 3340 351644 3352
rect 351696 3340 351702 3392
rect 354582 3340 354588 3392
rect 354640 3380 354646 3392
rect 472250 3380 472256 3392
rect 354640 3352 472256 3380
rect 354640 3340 354646 3352
rect 472250 3340 472256 3352
rect 472308 3340 472314 3392
rect 473354 3340 473360 3392
rect 473412 3380 473418 3392
rect 474550 3380 474556 3392
rect 473412 3352 474556 3380
rect 473412 3340 473418 3352
rect 474550 3340 474556 3352
rect 474608 3340 474614 3392
rect 481634 3340 481640 3392
rect 481692 3380 481698 3392
rect 482830 3380 482836 3392
rect 481692 3352 482836 3380
rect 481692 3340 481698 3352
rect 482830 3340 482836 3352
rect 482888 3340 482894 3392
rect 310606 3312 310612 3324
rect 306346 3284 310612 3312
rect 305365 3275 305423 3281
rect 310606 3272 310612 3284
rect 310664 3272 310670 3324
rect 311434 3272 311440 3324
rect 311492 3312 311498 3324
rect 313366 3312 313372 3324
rect 311492 3284 313372 3312
rect 311492 3272 311498 3284
rect 313366 3272 313372 3284
rect 313424 3272 313430 3324
rect 318702 3272 318708 3324
rect 318760 3312 318766 3324
rect 324501 3315 324559 3321
rect 324501 3312 324513 3315
rect 318760 3284 324513 3312
rect 318760 3272 318766 3284
rect 324501 3281 324513 3284
rect 324547 3281 324559 3315
rect 324501 3275 324559 3281
rect 329742 3272 329748 3324
rect 329800 3312 329806 3324
rect 334253 3315 334311 3321
rect 334253 3312 334265 3315
rect 329800 3284 334265 3312
rect 329800 3272 329806 3284
rect 334253 3281 334265 3284
rect 334299 3281 334311 3315
rect 334253 3275 334311 3281
rect 334345 3315 334403 3321
rect 334345 3281 334357 3315
rect 334391 3312 334403 3315
rect 362310 3312 362316 3324
rect 334391 3284 362316 3312
rect 334391 3281 334403 3284
rect 334345 3275 334403 3281
rect 362310 3272 362316 3284
rect 362368 3272 362374 3324
rect 398098 3272 398104 3324
rect 398156 3312 398162 3324
rect 514754 3312 514760 3324
rect 398156 3284 514760 3312
rect 398156 3272 398162 3284
rect 514754 3272 514760 3284
rect 514812 3272 514818 3324
rect 301516 3216 306374 3244
rect 301041 3207 301099 3213
rect 254302 3176 254308 3188
rect 71556 3148 92520 3176
rect 92584 3148 254308 3176
rect 71556 3136 71562 3148
rect 83274 3068 83280 3120
rect 83332 3108 83338 3120
rect 84102 3108 84108 3120
rect 83332 3080 84108 3108
rect 83332 3068 83338 3080
rect 84102 3068 84108 3080
rect 84160 3068 84166 3120
rect 78582 3000 78588 3052
rect 78640 3040 78646 3052
rect 92584 3040 92612 3148
rect 254302 3136 254308 3148
rect 254360 3136 254366 3188
rect 266538 3136 266544 3188
rect 266596 3176 266602 3188
rect 267642 3176 267648 3188
rect 266596 3148 267648 3176
rect 266596 3136 266602 3148
rect 267642 3136 267648 3148
rect 267700 3136 267706 3188
rect 285398 3136 285404 3188
rect 285456 3176 285462 3188
rect 299569 3179 299627 3185
rect 285456 3148 298140 3176
rect 285456 3136 285462 3148
rect 92750 3068 92756 3120
rect 92808 3108 92814 3120
rect 93762 3108 93768 3120
rect 92808 3080 93768 3108
rect 92808 3068 92814 3080
rect 93762 3068 93768 3080
rect 93820 3068 93826 3120
rect 93946 3068 93952 3120
rect 94004 3108 94010 3120
rect 95050 3108 95056 3120
rect 94004 3080 95056 3108
rect 94004 3068 94010 3080
rect 95050 3068 95056 3080
rect 95108 3068 95114 3120
rect 97442 3068 97448 3120
rect 97500 3108 97506 3120
rect 97902 3108 97908 3120
rect 97500 3080 97908 3108
rect 97500 3068 97506 3080
rect 97902 3068 97908 3080
rect 97960 3068 97966 3120
rect 98638 3068 98644 3120
rect 98696 3108 98702 3120
rect 99282 3108 99288 3120
rect 98696 3080 99288 3108
rect 98696 3068 98702 3080
rect 99282 3068 99288 3080
rect 99340 3068 99346 3120
rect 99834 3068 99840 3120
rect 99892 3108 99898 3120
rect 100662 3108 100668 3120
rect 99892 3080 100668 3108
rect 99892 3068 99898 3080
rect 100662 3068 100668 3080
rect 100720 3068 100726 3120
rect 256694 3108 256700 3120
rect 102060 3080 256700 3108
rect 102060 3040 102088 3080
rect 256694 3068 256700 3080
rect 256752 3068 256758 3120
rect 280706 3068 280712 3120
rect 280764 3108 280770 3120
rect 290645 3111 290703 3117
rect 290645 3108 290657 3111
rect 280764 3080 290657 3108
rect 280764 3068 280770 3080
rect 290645 3077 290657 3080
rect 290691 3077 290703 3111
rect 298005 3111 298063 3117
rect 298005 3108 298017 3111
rect 290645 3071 290703 3077
rect 290752 3080 298017 3108
rect 258442 3040 258448 3052
rect 78640 3012 92612 3040
rect 93826 3012 102088 3040
rect 102152 3012 258448 3040
rect 78640 3000 78646 3012
rect 89162 2932 89168 2984
rect 89220 2972 89226 2984
rect 93826 2972 93854 3012
rect 89220 2944 93854 2972
rect 89220 2932 89226 2944
rect 96246 2932 96252 2984
rect 96304 2972 96310 2984
rect 102152 2972 102180 3012
rect 258442 3000 258448 3012
rect 258500 3000 258506 3052
rect 290182 3000 290188 3052
rect 290240 3040 290246 3052
rect 290752 3040 290780 3080
rect 298005 3077 298017 3080
rect 298051 3077 298063 3111
rect 298112 3108 298140 3148
rect 299569 3145 299581 3179
rect 299615 3176 299627 3179
rect 305178 3176 305184 3188
rect 299615 3148 305184 3176
rect 299615 3145 299627 3148
rect 299569 3139 299627 3145
rect 305178 3136 305184 3148
rect 305236 3136 305242 3188
rect 306346 3176 306374 3216
rect 324038 3204 324044 3256
rect 324096 3244 324102 3256
rect 350442 3244 350448 3256
rect 324096 3216 350448 3244
rect 324096 3204 324102 3216
rect 350442 3204 350448 3216
rect 350500 3204 350506 3256
rect 353202 3204 353208 3256
rect 353260 3244 353266 3256
rect 465166 3244 465172 3256
rect 353260 3216 465172 3244
rect 353260 3204 353266 3216
rect 465166 3204 465172 3216
rect 465224 3204 465230 3256
rect 306466 3176 306472 3188
rect 306346 3148 306472 3176
rect 306466 3136 306472 3148
rect 306524 3136 306530 3188
rect 324130 3136 324136 3188
rect 324188 3176 324194 3188
rect 348050 3176 348056 3188
rect 324188 3148 348056 3176
rect 324188 3136 324194 3148
rect 348050 3136 348056 3148
rect 348108 3136 348114 3188
rect 351822 3136 351828 3188
rect 351880 3176 351886 3188
rect 458082 3176 458088 3188
rect 351880 3148 458088 3176
rect 351880 3136 351886 3148
rect 458082 3136 458088 3148
rect 458140 3136 458146 3188
rect 306558 3108 306564 3120
rect 298112 3080 306564 3108
rect 298005 3071 298063 3077
rect 306558 3068 306564 3080
rect 306616 3068 306622 3120
rect 318150 3068 318156 3120
rect 318208 3108 318214 3120
rect 320910 3108 320916 3120
rect 318208 3080 320916 3108
rect 318208 3068 318214 3080
rect 320910 3068 320916 3080
rect 320968 3068 320974 3120
rect 322842 3068 322848 3120
rect 322900 3108 322906 3120
rect 344554 3108 344560 3120
rect 322900 3080 344560 3108
rect 322900 3068 322906 3080
rect 344554 3068 344560 3080
rect 344612 3068 344618 3120
rect 347682 3068 347688 3120
rect 347740 3108 347746 3120
rect 443822 3108 443828 3120
rect 347740 3080 443828 3108
rect 347740 3068 347746 3080
rect 443822 3068 443828 3080
rect 443880 3068 443886 3120
rect 443914 3068 443920 3120
rect 443972 3108 443978 3120
rect 446493 3111 446551 3117
rect 443972 3080 446444 3108
rect 443972 3068 443978 3080
rect 290240 3012 290780 3040
rect 290240 3000 290246 3012
rect 293678 3000 293684 3052
rect 293736 3040 293742 3052
rect 309410 3040 309416 3052
rect 293736 3012 309416 3040
rect 293736 3000 293742 3012
rect 309410 3000 309416 3012
rect 309468 3000 309474 3052
rect 310238 3000 310244 3052
rect 310296 3040 310302 3052
rect 313458 3040 313464 3052
rect 310296 3012 313464 3040
rect 310296 3000 310302 3012
rect 313458 3000 313464 3012
rect 313516 3000 313522 3052
rect 322750 3000 322756 3052
rect 322808 3040 322814 3052
rect 343358 3040 343364 3052
rect 322808 3012 343364 3040
rect 322808 3000 322814 3012
rect 343358 3000 343364 3012
rect 343416 3000 343422 3052
rect 346302 3000 346308 3052
rect 346360 3040 346366 3052
rect 436738 3040 436744 3052
rect 346360 3012 436744 3040
rect 346360 3000 346366 3012
rect 436738 3000 436744 3012
rect 436796 3000 436802 3052
rect 436833 3043 436891 3049
rect 436833 3009 436845 3043
rect 436879 3040 436891 3043
rect 440421 3043 440479 3049
rect 440421 3040 440433 3043
rect 436879 3012 440433 3040
rect 436879 3009 436891 3012
rect 436833 3003 436891 3009
rect 440421 3009 440433 3012
rect 440467 3009 440479 3043
rect 440421 3003 440479 3009
rect 440878 3000 440884 3052
rect 440936 3040 440942 3052
rect 446309 3043 446367 3049
rect 446309 3040 446321 3043
rect 440936 3012 446321 3040
rect 440936 3000 440942 3012
rect 446309 3009 446321 3012
rect 446355 3009 446367 3043
rect 446416 3040 446444 3080
rect 446493 3077 446505 3111
rect 446539 3108 446551 3111
rect 454494 3108 454500 3120
rect 446539 3080 454500 3108
rect 446539 3077 446551 3080
rect 446493 3071 446551 3077
rect 454494 3068 454500 3080
rect 454552 3068 454558 3120
rect 446416 3012 447548 3040
rect 446309 3003 446367 3009
rect 96304 2944 102180 2972
rect 96304 2932 96310 2944
rect 102226 2932 102232 2984
rect 102284 2972 102290 2984
rect 103422 2972 103428 2984
rect 102284 2944 103428 2972
rect 102284 2932 102290 2944
rect 103422 2932 103428 2944
rect 103480 2932 103486 2984
rect 105722 2932 105728 2984
rect 105780 2972 105786 2984
rect 106182 2972 106188 2984
rect 105780 2944 106188 2972
rect 105780 2932 105786 2944
rect 106182 2932 106188 2944
rect 106240 2932 106246 2984
rect 106918 2932 106924 2984
rect 106976 2972 106982 2984
rect 107562 2972 107568 2984
rect 106976 2944 107568 2972
rect 106976 2932 106982 2944
rect 107562 2932 107568 2944
rect 107620 2932 107626 2984
rect 108114 2932 108120 2984
rect 108172 2972 108178 2984
rect 108942 2972 108948 2984
rect 108172 2944 108948 2972
rect 108172 2932 108178 2944
rect 108942 2932 108948 2944
rect 109000 2932 109006 2984
rect 109310 2932 109316 2984
rect 109368 2972 109374 2984
rect 110322 2972 110328 2984
rect 109368 2944 110328 2972
rect 109368 2932 109374 2944
rect 110322 2932 110328 2944
rect 110380 2932 110386 2984
rect 261110 2972 261116 2984
rect 110432 2944 261116 2972
rect 101030 2864 101036 2916
rect 101088 2904 101094 2916
rect 102042 2904 102048 2916
rect 101088 2876 102048 2904
rect 101088 2864 101094 2876
rect 102042 2864 102048 2876
rect 102100 2864 102106 2916
rect 103330 2864 103336 2916
rect 103388 2904 103394 2916
rect 110432 2904 110460 2944
rect 261110 2932 261116 2944
rect 261168 2932 261174 2984
rect 291378 2932 291384 2984
rect 291436 2972 291442 2984
rect 307846 2972 307852 2984
rect 291436 2944 307852 2972
rect 291436 2932 291442 2944
rect 307846 2932 307852 2944
rect 307904 2932 307910 2984
rect 321462 2932 321468 2984
rect 321520 2972 321526 2984
rect 340966 2972 340972 2984
rect 321520 2944 340972 2972
rect 321520 2932 321526 2944
rect 340966 2932 340972 2944
rect 341024 2932 341030 2984
rect 344922 2932 344928 2984
rect 344980 2972 344986 2984
rect 429654 2972 429660 2984
rect 344980 2944 429660 2972
rect 344980 2932 344986 2944
rect 429654 2932 429660 2944
rect 429712 2932 429718 2984
rect 429749 2975 429807 2981
rect 429749 2941 429761 2975
rect 429795 2972 429807 2975
rect 429795 2944 436784 2972
rect 429795 2941 429807 2944
rect 429749 2935 429807 2941
rect 103388 2876 110460 2904
rect 103388 2864 103394 2876
rect 110506 2864 110512 2916
rect 110564 2904 110570 2916
rect 262674 2904 262680 2916
rect 110564 2876 262680 2904
rect 110564 2864 110570 2876
rect 262674 2864 262680 2876
rect 262732 2864 262738 2916
rect 262950 2864 262956 2916
rect 263008 2904 263014 2916
rect 263502 2904 263508 2916
rect 263008 2876 263508 2904
rect 263008 2864 263014 2876
rect 263502 2864 263508 2876
rect 263560 2864 263566 2916
rect 294874 2864 294880 2916
rect 294932 2904 294938 2916
rect 309502 2904 309508 2916
rect 294932 2876 309508 2904
rect 294932 2864 294938 2876
rect 309502 2864 309508 2876
rect 309560 2864 309566 2916
rect 312630 2864 312636 2916
rect 312688 2904 312694 2916
rect 313550 2904 313556 2916
rect 312688 2876 313556 2904
rect 312688 2864 312694 2876
rect 313550 2864 313556 2876
rect 313608 2864 313614 2916
rect 317230 2864 317236 2916
rect 317288 2904 317294 2916
rect 324406 2904 324412 2916
rect 317288 2876 324412 2904
rect 317288 2864 317294 2876
rect 324406 2864 324412 2876
rect 324464 2864 324470 2916
rect 326890 2864 326896 2916
rect 326948 2904 326954 2916
rect 334345 2907 334403 2913
rect 334345 2904 334357 2907
rect 326948 2876 334357 2904
rect 326948 2864 326954 2876
rect 334345 2873 334357 2876
rect 334391 2873 334403 2907
rect 358722 2904 358728 2916
rect 334345 2867 334403 2873
rect 334452 2876 358728 2904
rect 114002 2796 114008 2848
rect 114060 2836 114066 2848
rect 114462 2836 114468 2848
rect 114060 2808 114468 2836
rect 114060 2796 114066 2808
rect 114462 2796 114468 2808
rect 114520 2796 114526 2848
rect 115198 2796 115204 2848
rect 115256 2836 115262 2848
rect 115842 2836 115848 2848
rect 115256 2808 115848 2836
rect 115256 2796 115262 2808
rect 115842 2796 115848 2808
rect 115900 2796 115906 2848
rect 116394 2796 116400 2848
rect 116452 2836 116458 2848
rect 117222 2836 117228 2848
rect 116452 2808 117228 2836
rect 116452 2796 116458 2808
rect 117222 2796 117228 2808
rect 117280 2796 117286 2848
rect 117590 2796 117596 2848
rect 117648 2836 117654 2848
rect 117648 2808 118740 2836
rect 117648 2796 117654 2808
rect 118712 2768 118740 2808
rect 118786 2796 118792 2848
rect 118844 2836 118850 2848
rect 119798 2836 119804 2848
rect 118844 2808 119804 2836
rect 118844 2796 118850 2808
rect 119798 2796 119804 2808
rect 119856 2796 119862 2848
rect 263870 2836 263876 2848
rect 119908 2808 263876 2836
rect 119908 2768 119936 2808
rect 263870 2796 263876 2808
rect 263928 2796 263934 2848
rect 292574 2796 292580 2848
rect 292632 2836 292638 2848
rect 298005 2839 298063 2845
rect 292632 2808 297956 2836
rect 292632 2796 292638 2808
rect 118712 2740 119936 2768
rect 297928 2768 297956 2808
rect 298005 2805 298017 2839
rect 298051 2836 298063 2839
rect 308214 2836 308220 2848
rect 298051 2808 308220 2836
rect 298051 2805 298063 2808
rect 298005 2799 298063 2805
rect 308214 2796 308220 2808
rect 308272 2796 308278 2848
rect 325602 2796 325608 2848
rect 325660 2836 325666 2848
rect 334253 2839 334311 2845
rect 334253 2836 334265 2839
rect 325660 2808 334265 2836
rect 325660 2796 325666 2808
rect 334253 2805 334265 2808
rect 334299 2805 334311 2839
rect 334253 2799 334311 2805
rect 301593 2771 301651 2777
rect 301593 2768 301605 2771
rect 297928 2740 301605 2768
rect 301593 2737 301605 2740
rect 301639 2737 301651 2771
rect 301593 2731 301651 2737
rect 333609 2771 333667 2777
rect 333609 2737 333621 2771
rect 333655 2768 333667 2771
rect 334452 2768 334480 2876
rect 358722 2864 358728 2876
rect 358780 2864 358786 2916
rect 383194 2864 383200 2916
rect 383252 2904 383258 2916
rect 408402 2904 408408 2916
rect 383252 2876 408408 2904
rect 383252 2864 383258 2876
rect 408402 2864 408408 2876
rect 408460 2864 408466 2916
rect 417418 2864 417424 2916
rect 417476 2904 417482 2916
rect 417476 2876 418752 2904
rect 417476 2864 417482 2876
rect 334529 2839 334587 2845
rect 334529 2805 334541 2839
rect 334575 2836 334587 2839
rect 355226 2836 355232 2848
rect 334575 2808 355232 2836
rect 334575 2805 334587 2808
rect 334529 2799 334587 2805
rect 355226 2796 355232 2808
rect 355284 2796 355290 2848
rect 405090 2796 405096 2848
rect 405148 2836 405154 2848
rect 418614 2836 418620 2848
rect 405148 2808 418620 2836
rect 405148 2796 405154 2808
rect 418614 2796 418620 2808
rect 418672 2796 418678 2848
rect 333655 2740 334480 2768
rect 418724 2768 418752 2876
rect 418798 2864 418804 2916
rect 418856 2904 418862 2916
rect 427081 2907 427139 2913
rect 427081 2904 427093 2907
rect 418856 2876 427093 2904
rect 418856 2864 418862 2876
rect 427081 2873 427093 2876
rect 427127 2873 427139 2907
rect 427081 2867 427139 2873
rect 427188 2876 432460 2904
rect 426989 2839 427047 2845
rect 426989 2836 427001 2839
rect 419092 2808 427001 2836
rect 419092 2768 419120 2808
rect 426989 2805 427001 2808
rect 427035 2805 427047 2839
rect 426989 2799 427047 2805
rect 418724 2740 419120 2768
rect 333655 2737 333667 2740
rect 333609 2731 333667 2737
rect 425790 2728 425796 2780
rect 425848 2768 425854 2780
rect 427188 2768 427216 2876
rect 427265 2839 427323 2845
rect 427265 2805 427277 2839
rect 427311 2836 427323 2839
rect 427311 2808 432368 2836
rect 427311 2805 427323 2808
rect 427265 2799 427323 2805
rect 425848 2740 427216 2768
rect 425848 2728 425854 2740
rect 432340 2700 432368 2808
rect 432432 2768 432460 2876
rect 432506 2864 432512 2916
rect 432564 2904 432570 2916
rect 433242 2904 433248 2916
rect 432564 2876 433248 2904
rect 432564 2864 432570 2876
rect 433242 2864 433248 2876
rect 433300 2864 433306 2916
rect 436649 2907 436707 2913
rect 436649 2904 436661 2907
rect 433352 2876 436661 2904
rect 433352 2768 433380 2876
rect 436649 2873 436661 2876
rect 436695 2873 436707 2907
rect 436756 2904 436784 2944
rect 436922 2932 436928 2984
rect 436980 2972 436986 2984
rect 447410 2972 447416 2984
rect 436980 2944 447416 2972
rect 436980 2932 436986 2944
rect 447410 2932 447416 2944
rect 447468 2932 447474 2984
rect 447520 2972 447548 3012
rect 447778 3000 447784 3052
rect 447836 3040 447842 3052
rect 468662 3040 468668 3052
rect 447836 3012 468668 3040
rect 447836 3000 447842 3012
rect 468662 3000 468668 3012
rect 468720 3000 468726 3052
rect 461578 2972 461584 2984
rect 447520 2944 461584 2972
rect 461578 2932 461584 2944
rect 461636 2932 461642 2984
rect 479334 2904 479340 2916
rect 436756 2876 479340 2904
rect 436649 2867 436707 2873
rect 479334 2864 479340 2876
rect 479392 2864 479398 2916
rect 450906 2836 450912 2848
rect 432432 2740 433380 2768
rect 433444 2808 450912 2836
rect 433444 2700 433472 2808
rect 450906 2796 450912 2808
rect 450964 2796 450970 2848
rect 450998 2796 451004 2848
rect 451056 2836 451062 2848
rect 475746 2836 475752 2848
rect 451056 2808 475752 2836
rect 451056 2796 451062 2808
rect 475746 2796 475752 2808
rect 475804 2796 475810 2848
rect 432340 2672 433472 2700
<< via1 >>
rect 170312 700952 170364 701004
rect 316040 700952 316092 701004
rect 154120 700884 154172 700936
rect 312544 700884 312596 700936
rect 299388 700816 299440 700868
rect 462320 700816 462372 700868
rect 300768 700748 300820 700800
rect 478512 700748 478564 700800
rect 137836 700680 137888 700732
rect 317420 700680 317472 700732
rect 298008 700612 298060 700664
rect 494796 700612 494848 700664
rect 105452 700544 105504 700596
rect 320180 700544 320232 700596
rect 89168 700476 89220 700528
rect 315304 700476 315356 700528
rect 295248 700408 295300 700460
rect 527180 700408 527232 700460
rect 296628 700340 296680 700392
rect 543464 700340 543516 700392
rect 72976 700272 73028 700324
rect 321560 700272 321612 700324
rect 302148 700204 302200 700256
rect 429844 700204 429896 700256
rect 202788 700136 202840 700188
rect 313280 700136 313332 700188
rect 304908 700068 304960 700120
rect 413652 700068 413704 700120
rect 303528 700000 303580 700052
rect 397460 700000 397512 700052
rect 235172 699932 235224 699984
rect 311992 699932 312044 699984
rect 306288 699864 306340 699916
rect 364984 699864 365036 699916
rect 267648 699796 267700 699848
rect 310520 699796 310572 699848
rect 307668 699728 307720 699780
rect 332508 699728 332560 699780
rect 300124 699660 300176 699712
rect 309140 699660 309192 699712
rect 292488 696940 292540 696992
rect 580172 696940 580224 696992
rect 292396 683204 292448 683256
rect 580172 683204 580224 683256
rect 3424 683136 3476 683188
rect 328460 683136 328512 683188
rect 291108 670760 291160 670812
rect 580172 670760 580224 670812
rect 3516 670692 3568 670744
rect 323584 670692 323636 670744
rect 3424 656888 3476 656940
rect 329840 656888 329892 656940
rect 288348 643084 288400 643136
rect 580172 643084 580224 643136
rect 3424 632068 3476 632120
rect 332600 632068 332652 632120
rect 289728 630640 289780 630692
rect 580172 630640 580224 630692
rect 3148 618264 3200 618316
rect 327724 618264 327776 618316
rect 286968 616836 287020 616888
rect 580172 616836 580224 616888
rect 3240 605820 3292 605872
rect 332692 605820 332744 605872
rect 284116 590656 284168 590708
rect 579804 590656 579856 590708
rect 3332 579640 3384 579692
rect 335360 579640 335412 579692
rect 285588 576852 285640 576904
rect 580172 576852 580224 576904
rect 3424 565836 3476 565888
rect 331864 565836 331916 565888
rect 282828 563048 282880 563100
rect 579804 563048 579856 563100
rect 3424 553392 3476 553444
rect 336740 553392 336792 553444
rect 280068 536800 280120 536852
rect 580172 536800 580224 536852
rect 3424 527144 3476 527196
rect 339500 527144 339552 527196
rect 281448 524424 281500 524476
rect 580172 524424 580224 524476
rect 3424 514768 3476 514820
rect 334624 514768 334676 514820
rect 278688 510620 278740 510672
rect 580172 510620 580224 510672
rect 3056 500964 3108 501016
rect 340880 500964 340932 501016
rect 285128 491240 285180 491292
rect 285588 491240 285640 491292
rect 286416 491240 286468 491292
rect 286968 491240 287020 491292
rect 287704 491240 287756 491292
rect 288348 491240 288400 491292
rect 288992 491240 289044 491292
rect 289728 491240 289780 491292
rect 290280 491240 290332 491292
rect 291108 491240 291160 491292
rect 291568 491240 291620 491292
rect 292488 491240 292540 491292
rect 305828 491240 305880 491292
rect 306288 491240 306340 491292
rect 307116 491240 307168 491292
rect 307668 491240 307720 491292
rect 327724 491240 327776 491292
rect 334900 491240 334952 491292
rect 284208 491172 284260 491224
rect 311900 491172 311952 491224
rect 312544 491172 312596 491224
rect 319352 491172 319404 491224
rect 319444 491172 319496 491224
rect 327172 491172 327224 491224
rect 331864 491172 331916 491224
rect 338764 491172 338816 491224
rect 308404 491104 308456 491156
rect 347780 491104 347832 491156
rect 219348 491036 219400 491088
rect 315212 491036 315264 491088
rect 315304 491036 315356 491088
rect 323308 491036 323360 491088
rect 323584 491036 323636 491088
rect 331220 491036 331272 491088
rect 334624 491036 334676 491088
rect 342720 491036 342772 491088
rect 273168 490968 273220 491020
rect 385960 490968 386012 491020
rect 271788 490900 271840 490952
rect 386052 490900 386104 490952
rect 7932 490832 7984 490884
rect 346584 490832 346636 490884
rect 5448 490764 5500 490816
rect 347964 490764 348016 490816
rect 5356 490696 5408 490748
rect 349160 490696 349212 490748
rect 5264 490628 5316 490680
rect 351920 490628 351972 490680
rect 3332 490560 3384 490612
rect 350540 490560 350592 490612
rect 4068 490492 4120 490544
rect 354312 490492 354364 490544
rect 3976 490424 4028 490476
rect 353300 490424 353352 490476
rect 6552 490356 6604 490408
rect 356888 490356 356940 490408
rect 3884 490288 3936 490340
rect 358176 490288 358228 490340
rect 6460 490220 6512 490272
rect 360752 490220 360804 490272
rect 3792 490152 3844 490204
rect 362132 490152 362184 490204
rect 6368 490084 6420 490136
rect 364708 490084 364760 490136
rect 3608 490016 3660 490068
rect 365996 490016 366048 490068
rect 6276 489948 6328 490000
rect 368572 489948 368624 490000
rect 3424 489880 3476 489932
rect 369860 489880 369912 489932
rect 275928 488452 275980 488504
rect 384120 488452 384172 488504
rect 274548 488384 274600 488436
rect 383200 488384 383252 488436
rect 277124 488316 277176 488368
rect 386144 488316 386196 488368
rect 268292 488248 268344 488300
rect 385868 488248 385920 488300
rect 255228 488180 255280 488232
rect 383384 488180 383436 488232
rect 247592 488112 247644 488164
rect 383108 488112 383160 488164
rect 248880 488044 248932 488096
rect 384672 488044 384724 488096
rect 243728 487976 243780 488028
rect 383016 487976 383068 488028
rect 245016 487908 245068 487960
rect 384580 487908 384632 487960
rect 239864 487840 239916 487892
rect 382924 487840 382976 487892
rect 235908 487772 235960 487824
rect 393964 487772 394016 487824
rect 269258 487704 269310 487756
rect 580908 487704 580960 487756
rect 250168 487636 250220 487688
rect 580356 487636 580408 487688
rect 4712 487568 4764 487620
rect 344008 487568 344060 487620
rect 345296 487611 345348 487620
rect 345296 487577 345305 487611
rect 345305 487577 345339 487611
rect 345339 487577 345348 487611
rect 345296 487568 345348 487577
rect 4988 487500 5040 487552
rect 371240 487568 371292 487620
rect 355600 487543 355652 487552
rect 355600 487509 355609 487543
rect 355609 487509 355643 487543
rect 355643 487509 355652 487543
rect 355600 487500 355652 487509
rect 359464 487543 359516 487552
rect 359464 487509 359473 487543
rect 359473 487509 359507 487543
rect 359507 487509 359516 487543
rect 359464 487500 359516 487509
rect 363420 487543 363472 487552
rect 363420 487509 363429 487543
rect 363429 487509 363463 487543
rect 363463 487509 363472 487543
rect 363420 487500 363472 487509
rect 367284 487543 367336 487552
rect 367284 487509 367293 487543
rect 367293 487509 367327 487543
rect 367327 487509 367336 487543
rect 367284 487500 367336 487509
rect 7748 487432 7800 487484
rect 376300 487500 376352 487552
rect 4896 487364 4948 487416
rect 375012 487364 375064 487416
rect 7564 487296 7616 487348
rect 380164 487296 380216 487348
rect 7656 487228 7708 487280
rect 381452 487228 381504 487280
rect 4804 487160 4856 487212
rect 378876 487160 378928 487212
rect 270868 487092 270920 487144
rect 384212 487092 384264 487144
rect 241152 487024 241204 487076
rect 257896 487067 257948 487076
rect 246304 486956 246356 487008
rect 257896 487033 257905 487067
rect 257905 487033 257939 487067
rect 257939 487033 257948 487067
rect 257896 487024 257948 487033
rect 259276 487024 259328 487076
rect 251272 486956 251324 487008
rect 252560 486999 252612 487008
rect 252560 486965 252569 486999
rect 252569 486965 252603 486999
rect 252603 486965 252612 486999
rect 252560 486956 252612 486965
rect 253848 486999 253900 487008
rect 253848 486965 253857 486999
rect 253857 486965 253891 486999
rect 253891 486965 253900 486999
rect 253848 486956 253900 486965
rect 256608 486956 256660 487008
rect 260564 486956 260616 487008
rect 261852 486999 261904 487008
rect 261852 486965 261861 486999
rect 261861 486965 261895 486999
rect 261895 486965 261904 486999
rect 261852 486956 261904 486965
rect 263140 487024 263192 487076
rect 264428 486999 264480 487008
rect 264428 486965 264437 486999
rect 264437 486965 264471 486999
rect 264471 486965 264480 486999
rect 264428 486956 264480 486965
rect 265716 486999 265768 487008
rect 265716 486965 265725 486999
rect 265725 486965 265759 486999
rect 265759 486965 265768 486999
rect 265716 486956 265768 486965
rect 267004 487024 267056 487076
rect 384948 487024 385000 487076
rect 383568 486956 383620 487008
rect 383476 486888 383528 486940
rect 385776 486820 385828 486872
rect 384856 486752 384908 486804
rect 383292 486684 383344 486736
rect 384764 486616 384816 486668
rect 384396 486548 384448 486600
rect 580724 486480 580776 486532
rect 580816 486412 580868 486464
rect 580632 486344 580684 486396
rect 580540 486276 580592 486328
rect 580448 486208 580500 486260
rect 580264 486140 580316 486192
rect 6644 486072 6696 486124
rect 5172 486004 5224 486056
rect 5080 485936 5132 485988
rect 3700 485868 3752 485920
rect 3516 485800 3568 485852
rect 384120 485732 384172 485784
rect 580172 485732 580224 485784
rect 2780 475668 2832 475720
rect 4712 475668 4764 475720
rect 386144 471928 386196 471980
rect 580172 471928 580224 471980
rect 3240 462680 3292 462732
rect 7932 462680 7984 462732
rect 383200 458124 383252 458176
rect 580172 458124 580224 458176
rect 3240 449556 3292 449608
rect 6644 449556 6696 449608
rect 386052 431876 386104 431928
rect 580172 431876 580224 431928
rect 2780 423580 2832 423632
rect 5448 423580 5500 423632
rect 385960 419432 386012 419484
rect 580172 419432 580224 419484
rect 384212 405628 384264 405680
rect 580172 405628 580224 405680
rect 2780 397536 2832 397588
rect 5356 397536 5408 397588
rect 385868 379448 385920 379500
rect 579988 379448 580040 379500
rect 2780 371424 2832 371476
rect 5264 371424 5316 371476
rect 384948 353200 385000 353252
rect 580172 353200 580224 353252
rect 251226 337764 251278 337816
rect 251548 337764 251600 337816
rect 265026 337764 265078 337816
rect 265256 337764 265308 337816
rect 75828 336676 75880 336728
rect 284300 336744 284352 336796
rect 284668 336744 284720 336796
rect 293960 336744 294012 336796
rect 294788 336744 294840 336796
rect 337936 336744 337988 336796
rect 376116 336744 376168 336796
rect 253756 336676 253808 336728
rect 258172 336676 258224 336728
rect 258540 336676 258592 336728
rect 68928 336608 68980 336660
rect 252008 336608 252060 336660
rect 278320 336676 278372 336728
rect 281540 336676 281592 336728
rect 281908 336676 281960 336728
rect 282276 336676 282328 336728
rect 305184 336676 305236 336728
rect 313372 336676 313424 336728
rect 313556 336676 313608 336728
rect 317788 336676 317840 336728
rect 320824 336676 320876 336728
rect 321192 336676 321244 336728
rect 321468 336676 321520 336728
rect 322020 336676 322072 336728
rect 322756 336676 322808 336728
rect 323860 336676 323912 336728
rect 324228 336676 324280 336728
rect 325240 336676 325292 336728
rect 325516 336676 325568 336728
rect 327632 336676 327684 336728
rect 328276 336676 328328 336728
rect 329472 336676 329524 336728
rect 329748 336676 329800 336728
rect 330668 336676 330720 336728
rect 330852 336676 330904 336728
rect 331864 336676 331916 336728
rect 332324 336676 332376 336728
rect 334900 336676 334952 336728
rect 335268 336676 335320 336728
rect 337660 336676 337712 336728
rect 338764 336676 338816 336728
rect 339132 336676 339184 336728
rect 339224 336676 339276 336728
rect 339408 336676 339460 336728
rect 340512 336676 340564 336728
rect 340788 336676 340840 336728
rect 341432 336676 341484 336728
rect 342168 336676 342220 336728
rect 342628 336676 342680 336728
rect 343364 336676 343416 336728
rect 62028 336540 62080 336592
rect 250168 336540 250220 336592
rect 53748 336472 53800 336524
rect 248420 336472 248472 336524
rect 267648 336608 267700 336660
rect 302240 336608 302292 336660
rect 318800 336608 318852 336660
rect 322204 336608 322256 336660
rect 324688 336608 324740 336660
rect 325332 336608 325384 336660
rect 326436 336608 326488 336660
rect 326804 336608 326856 336660
rect 328828 336608 328880 336660
rect 329656 336608 329708 336660
rect 330024 336608 330076 336660
rect 330944 336608 330996 336660
rect 331956 336608 332008 336660
rect 332508 336608 332560 336660
rect 334256 336608 334308 336660
rect 335084 336608 335136 336660
rect 339960 336608 340012 336660
rect 340696 336608 340748 336660
rect 342904 336608 342956 336660
rect 343548 336608 343600 336660
rect 263508 336540 263560 336592
rect 301320 336540 301372 336592
rect 311164 336540 311216 336592
rect 311900 336540 311952 336592
rect 318064 336540 318116 336592
rect 318616 336540 318668 336592
rect 324964 336540 325016 336592
rect 325608 336540 325660 336592
rect 325884 336540 325936 336592
rect 326988 336540 327040 336592
rect 337568 336540 337620 336592
rect 338764 336540 338816 336592
rect 341156 336540 341208 336592
rect 405096 336676 405148 336728
rect 343824 336608 343876 336660
rect 344928 336608 344980 336660
rect 345296 336608 345348 336660
rect 346032 336608 346084 336660
rect 346860 336608 346912 336660
rect 347504 336608 347556 336660
rect 348608 336608 348660 336660
rect 349068 336608 349120 336660
rect 349804 336608 349856 336660
rect 350264 336608 350316 336660
rect 351276 336608 351328 336660
rect 351736 336608 351788 336660
rect 352932 336608 352984 336660
rect 353116 336608 353168 336660
rect 354036 336608 354088 336660
rect 354496 336608 354548 336660
rect 345940 336540 345992 336592
rect 346216 336540 346268 336592
rect 347412 336540 347464 336592
rect 347688 336540 347740 336592
rect 348056 336540 348108 336592
rect 348884 336540 348936 336592
rect 349528 336540 349580 336592
rect 350448 336540 350500 336592
rect 350724 336540 350776 336592
rect 351552 336540 351604 336592
rect 417424 336608 417476 336660
rect 354864 336540 354916 336592
rect 355692 336540 355744 336592
rect 359648 336540 359700 336592
rect 360108 336540 360160 336592
rect 360568 336540 360620 336592
rect 361304 336540 361356 336592
rect 362408 336540 362460 336592
rect 362684 336540 362736 336592
rect 363236 336540 363288 336592
rect 364156 336540 364208 336592
rect 425704 336540 425756 336592
rect 42708 336404 42760 336456
rect 245384 336404 245436 336456
rect 37188 336336 37240 336388
rect 243912 336336 243964 336388
rect 245016 336336 245068 336388
rect 300400 336472 300452 336524
rect 307668 336472 307720 336524
rect 312360 336472 312412 336524
rect 316592 336472 316644 336524
rect 320916 336472 320968 336524
rect 341984 336472 342036 336524
rect 416044 336472 416096 336524
rect 254584 336404 254636 336456
rect 296812 336404 296864 336456
rect 316868 336404 316920 336456
rect 322388 336404 322440 336456
rect 344744 336404 344796 336456
rect 429844 336404 429896 336456
rect 256608 336336 256660 336388
rect 299572 336336 299624 336388
rect 319996 336336 320048 336388
rect 335728 336336 335780 336388
rect 345664 336336 345716 336388
rect 346308 336336 346360 336388
rect 351000 336336 351052 336388
rect 351828 336336 351880 336388
rect 432604 336336 432656 336388
rect 44088 336268 44140 336320
rect 245660 336268 245712 336320
rect 246396 336268 246448 336320
rect 290280 336268 290332 336320
rect 315396 336268 315448 336320
rect 316316 336268 316368 336320
rect 319904 336268 319956 336320
rect 334440 336268 334492 336320
rect 344100 336268 344152 336320
rect 344744 336268 344796 336320
rect 349160 336268 349212 336320
rect 352840 336268 352892 336320
rect 353208 336268 353260 336320
rect 436744 336268 436796 336320
rect 35808 336200 35860 336252
rect 243636 336200 243688 336252
rect 251824 336200 251876 336252
rect 295984 336200 296036 336252
rect 319260 336200 319312 336252
rect 324964 336200 325016 336252
rect 350080 336200 350132 336252
rect 440884 336200 440936 336252
rect 28908 336132 28960 336184
rect 241796 336132 241848 336184
rect 244924 336132 244976 336184
rect 290096 336132 290148 336184
rect 320732 336132 320784 336184
rect 338580 336132 338632 336184
rect 346400 336132 346452 336184
rect 351920 336132 351972 336184
rect 443644 336132 443696 336184
rect 19248 336064 19300 336116
rect 239404 336064 239456 336116
rect 252468 336064 252520 336116
rect 298652 336064 298704 336116
rect 315948 336064 316000 336116
rect 318892 336064 318944 336116
rect 321100 336064 321152 336116
rect 339868 336064 339920 336116
rect 348332 336064 348384 336116
rect 353668 336064 353720 336116
rect 447784 336064 447836 336116
rect 20628 335996 20680 336048
rect 240140 335996 240192 336048
rect 249064 335996 249116 336048
rect 296536 335996 296588 336048
rect 303528 335996 303580 336048
rect 311532 335996 311584 336048
rect 316132 335996 316184 336048
rect 317972 335996 318024 336048
rect 322848 335996 322900 336048
rect 346768 335996 346820 336048
rect 357900 335996 357952 336048
rect 358728 335996 358780 336048
rect 359096 335996 359148 336048
rect 359924 335996 359976 336048
rect 361764 335996 361816 336048
rect 362592 335996 362644 336048
rect 450544 335996 450596 336048
rect 82728 335928 82780 335980
rect 255596 335928 255648 335980
rect 260748 335928 260800 335980
rect 269028 335928 269080 335980
rect 302792 335928 302844 335980
rect 323216 335928 323268 335980
rect 324136 335928 324188 335980
rect 337292 335928 337344 335980
rect 337752 335928 337804 335980
rect 343180 335928 343232 335980
rect 343456 335928 343508 335980
rect 93768 335860 93820 335912
rect 258356 335860 258408 335912
rect 271236 335860 271288 335912
rect 301964 335860 302016 335912
rect 340236 335860 340288 335912
rect 391204 335928 391256 335980
rect 86868 335792 86920 335844
rect 256424 335792 256476 335844
rect 274548 335792 274600 335844
rect 303988 335792 304040 335844
rect 327356 335792 327408 335844
rect 328092 335792 328144 335844
rect 333060 335792 333112 335844
rect 333888 335792 333940 335844
rect 338488 335792 338540 335844
rect 362040 335792 362092 335844
rect 362868 335792 362920 335844
rect 364248 335792 364300 335844
rect 366272 335792 366324 335844
rect 366732 335792 366784 335844
rect 366916 335792 366968 335844
rect 100668 335724 100720 335776
rect 260012 335724 260064 335776
rect 285588 335724 285640 335776
rect 306748 335724 306800 335776
rect 335544 335724 335596 335776
rect 336556 335724 336608 335776
rect 356428 335724 356480 335776
rect 107568 335656 107620 335708
rect 261852 335656 261904 335708
rect 288348 335656 288400 335708
rect 307760 335656 307812 335708
rect 330392 335656 330444 335708
rect 331128 335656 331180 335708
rect 331588 335656 331640 335708
rect 332232 335656 332284 335708
rect 336924 335656 336976 335708
rect 337936 335656 337988 335708
rect 355232 335656 355284 335708
rect 355876 335656 355928 335708
rect 361212 335656 361264 335708
rect 361488 335656 361540 335708
rect 114468 335588 114520 335640
rect 263600 335588 263652 335640
rect 286968 335588 287020 335640
rect 307300 335588 307352 335640
rect 315120 335588 315172 335640
rect 316132 335588 316184 335640
rect 355508 335588 355560 335640
rect 121368 335520 121420 335572
rect 265440 335520 265492 335572
rect 289728 335520 289780 335572
rect 307944 335520 307996 335572
rect 319628 335520 319680 335572
rect 320088 335520 320140 335572
rect 366548 335724 366600 335776
rect 367008 335724 367060 335776
rect 365996 335656 366048 335708
rect 366916 335656 366968 335708
rect 367744 335792 367796 335844
rect 368204 335792 368256 335844
rect 369216 335792 369268 335844
rect 369676 335792 369728 335844
rect 370780 335792 370832 335844
rect 367468 335724 367520 335776
rect 368296 335724 368348 335776
rect 368664 335724 368716 335776
rect 369492 335724 369544 335776
rect 372528 335724 372580 335776
rect 378784 335724 378836 335776
rect 379244 335724 379296 335776
rect 380348 335860 380400 335912
rect 380624 335860 380676 335912
rect 379980 335792 380032 335844
rect 380808 335792 380860 335844
rect 381176 335860 381228 335912
rect 382096 335860 382148 335912
rect 383200 335792 383252 335844
rect 411904 335792 411956 335844
rect 413284 335724 413336 335776
rect 405004 335656 405056 335708
rect 364800 335588 364852 335640
rect 365536 335588 365588 335640
rect 368940 335588 368992 335640
rect 193864 335452 193916 335504
rect 266360 335452 266412 335504
rect 322296 335452 322348 335504
rect 322848 335452 322900 335504
rect 191104 335384 191156 335436
rect 265992 335384 266044 335436
rect 318984 335384 319036 335436
rect 327724 335452 327776 335504
rect 363880 335452 363932 335504
rect 364248 335452 364300 335504
rect 326528 335384 326580 335436
rect 326896 335384 326948 335436
rect 336096 335384 336148 335436
rect 336464 335384 336516 335436
rect 243544 335316 243596 335368
rect 277400 335316 277452 335368
rect 315672 335316 315724 335368
rect 317512 335316 317564 335368
rect 352196 335316 352248 335368
rect 365352 335520 365404 335572
rect 398104 335588 398156 335640
rect 377404 335520 377456 335572
rect 403624 335520 403676 335572
rect 399484 335452 399536 335504
rect 371976 335384 372028 335436
rect 372528 335384 372580 335436
rect 372804 335384 372856 335436
rect 373908 335384 373960 335436
rect 377036 335384 377088 335436
rect 370412 335316 370464 335368
rect 370872 335316 370924 335368
rect 370964 335316 371016 335368
rect 371148 335316 371200 335368
rect 371608 335316 371660 335368
rect 372160 335316 372212 335368
rect 373172 335316 373224 335368
rect 373540 335316 373592 335368
rect 373632 335316 373684 335368
rect 373816 335316 373868 335368
rect 374644 335316 374696 335368
rect 375012 335316 375064 335368
rect 375104 335316 375156 335368
rect 375288 335316 375340 335368
rect 375840 335316 375892 335368
rect 376484 335316 376536 335368
rect 377312 335316 377364 335368
rect 378048 335316 378100 335368
rect 378508 335384 378560 335436
rect 379244 335384 379296 335436
rect 396724 335384 396776 335436
rect 379060 335316 379112 335368
rect 379336 335316 379388 335368
rect 353116 335180 353168 335232
rect 261116 330760 261168 330812
rect 272156 330760 272208 330812
rect 332416 330624 332468 330676
rect 261116 330556 261168 330608
rect 272156 330556 272208 330608
rect 309140 330556 309192 330608
rect 310336 330556 310388 330608
rect 254124 330488 254176 330540
rect 254952 330488 255004 330540
rect 256700 330488 256752 330540
rect 257344 330488 257396 330540
rect 259736 330488 259788 330540
rect 260656 330488 260708 330540
rect 261024 330488 261076 330540
rect 261576 330488 261628 330540
rect 262496 330488 262548 330540
rect 263324 330488 263376 330540
rect 265072 330488 265124 330540
rect 265716 330488 265768 330540
rect 266452 330488 266504 330540
rect 266912 330488 266964 330540
rect 267924 330488 267976 330540
rect 268752 330488 268804 330540
rect 269120 330488 269172 330540
rect 269580 330488 269632 330540
rect 270776 330488 270828 330540
rect 271696 330488 271748 330540
rect 272064 330488 272116 330540
rect 272616 330488 272668 330540
rect 302424 330488 302476 330540
rect 303436 330488 303488 330540
rect 305184 330488 305236 330540
rect 305828 330488 305880 330540
rect 307852 330488 307904 330540
rect 308496 330488 308548 330540
rect 309232 330488 309284 330540
rect 309692 330488 309744 330540
rect 313280 330488 313332 330540
rect 314200 330488 314252 330540
rect 266544 330420 266596 330472
rect 267188 330420 267240 330472
rect 267740 330420 267792 330472
rect 268384 330420 268436 330472
rect 269212 330420 269264 330472
rect 269948 330420 270000 330472
rect 270592 330420 270644 330472
rect 271420 330420 271472 330472
rect 271880 330420 271932 330472
rect 272892 330420 272944 330472
rect 307944 330420 307996 330472
rect 308772 330420 308824 330472
rect 309324 330420 309376 330472
rect 309968 330420 310020 330472
rect 320456 330420 320508 330472
rect 321376 330420 321428 330472
rect 323768 330420 323820 330472
rect 324044 330420 324096 330472
rect 326160 330420 326212 330472
rect 326712 330420 326764 330472
rect 332232 330420 332284 330472
rect 370136 330488 370188 330540
rect 371056 330488 371108 330540
rect 374368 330488 374420 330540
rect 375196 330488 375248 330540
rect 376392 330488 376444 330540
rect 376668 330488 376720 330540
rect 357164 330420 357216 330472
rect 357440 330420 357492 330472
rect 302332 328924 302384 328976
rect 303160 328924 303212 328976
rect 255412 327632 255464 327684
rect 256148 327632 256200 327684
rect 288716 326816 288768 326868
rect 256884 326748 256936 326800
rect 257620 326748 257672 326800
rect 278780 326680 278832 326732
rect 279056 326680 279108 326732
rect 284484 326680 284536 326732
rect 284760 326680 284812 326732
rect 293868 326680 293920 326732
rect 294420 326680 294472 326732
rect 288716 326612 288768 326664
rect 262404 326544 262456 326596
rect 263048 326544 263100 326596
rect 287060 326476 287112 326528
rect 287336 326476 287388 326528
rect 294052 326476 294104 326528
rect 294328 326476 294380 326528
rect 295524 326519 295576 326528
rect 295524 326485 295533 326519
rect 295533 326485 295567 326519
rect 295567 326485 295576 326519
rect 295524 326476 295576 326485
rect 244556 326408 244608 326460
rect 245108 326408 245160 326460
rect 245936 326408 245988 326460
rect 246580 326408 246632 326460
rect 247316 326408 247368 326460
rect 248052 326408 248104 326460
rect 252744 326408 252796 326460
rect 253480 326408 253532 326460
rect 276204 326408 276256 326460
rect 277124 326408 277176 326460
rect 280252 326408 280304 326460
rect 280988 326408 281040 326460
rect 281724 326408 281776 326460
rect 282460 326408 282512 326460
rect 283104 326408 283156 326460
rect 283932 326408 283984 326460
rect 284392 326408 284444 326460
rect 285496 326408 285548 326460
rect 288440 326408 288492 326460
rect 289084 326408 289136 326460
rect 291200 326408 291252 326460
rect 291752 326408 291804 326460
rect 296904 326408 296956 326460
rect 297732 326408 297784 326460
rect 234712 326340 234764 326392
rect 235540 326340 235592 326392
rect 236092 326340 236144 326392
rect 236736 326340 236788 326392
rect 237380 326340 237432 326392
rect 238484 326340 238536 326392
rect 238852 326340 238904 326392
rect 239680 326340 239732 326392
rect 240324 326340 240376 326392
rect 240876 326340 240928 326392
rect 241612 326340 241664 326392
rect 242072 326340 242124 326392
rect 244372 326340 244424 326392
rect 244832 326340 244884 326392
rect 245752 326340 245804 326392
rect 246304 326340 246356 326392
rect 247224 326340 247276 326392
rect 247776 326340 247828 326392
rect 248512 326340 248564 326392
rect 249616 326340 249668 326392
rect 249892 326340 249944 326392
rect 250812 326340 250864 326392
rect 251272 326340 251324 326392
rect 252284 326340 252336 326392
rect 252652 326340 252704 326392
rect 253204 326340 253256 326392
rect 273444 326340 273496 326392
rect 274088 326340 274140 326392
rect 276112 326340 276164 326392
rect 276756 326340 276808 326392
rect 278872 326340 278924 326392
rect 279516 326340 279568 326392
rect 280436 326340 280488 326392
rect 281264 326340 281316 326392
rect 281632 326340 281684 326392
rect 282184 326340 282236 326392
rect 283012 326340 283064 326392
rect 283656 326340 283708 326392
rect 284576 326340 284628 326392
rect 285220 326340 285272 326392
rect 287336 326340 287388 326392
rect 287888 326340 287940 326392
rect 288624 326340 288676 326392
rect 289360 326340 289412 326392
rect 289912 326340 289964 326392
rect 290556 326340 290608 326392
rect 291476 326340 291528 326392
rect 292396 326340 292448 326392
rect 296812 326340 296864 326392
rect 297456 326340 297508 326392
rect 298284 326340 298336 326392
rect 299204 326340 299256 326392
rect 299572 326340 299624 326392
rect 300124 326340 300176 326392
rect 247040 326272 247092 326324
rect 247500 326272 247552 326324
rect 291292 326272 291344 326324
rect 292028 326272 292080 326324
rect 292580 324232 292632 324284
rect 293592 324232 293644 324284
rect 242992 323552 243044 323604
rect 243176 323552 243228 323604
rect 285680 323552 285732 323604
rect 286416 323552 286468 323604
rect 288532 323552 288584 323604
rect 288808 323552 288860 323604
rect 295524 323595 295576 323604
rect 295524 323561 295533 323595
rect 295533 323561 295567 323595
rect 295567 323561 295576 323595
rect 295524 323552 295576 323561
rect 273260 323280 273312 323332
rect 273812 323280 273864 323332
rect 236184 323144 236236 323196
rect 237012 323144 237064 323196
rect 240232 321852 240284 321904
rect 240600 321852 240652 321904
rect 287152 321784 287204 321836
rect 288164 321784 288216 321836
rect 251456 320696 251508 320748
rect 251640 320696 251692 320748
rect 2780 319812 2832 319864
rect 5172 319812 5224 319864
rect 238944 319540 238996 319592
rect 239128 319540 239180 319592
rect 383568 299412 383620 299464
rect 580172 299412 580224 299464
rect 3148 293768 3200 293820
rect 6552 293768 6604 293820
rect 385776 273164 385828 273216
rect 580172 273164 580224 273216
rect 2780 267248 2832 267300
rect 5080 267248 5132 267300
rect 383476 245556 383528 245608
rect 580172 245556 580224 245608
rect 3240 241068 3292 241120
rect 6460 241068 6512 241120
rect 384856 233180 384908 233232
rect 579988 233180 580040 233232
rect 383384 206932 383436 206984
rect 580172 206932 580224 206984
rect 384764 193128 384816 193180
rect 580172 193128 580224 193180
rect 3240 188844 3292 188896
rect 6368 188844 6420 188896
rect 383292 166948 383344 167000
rect 580172 166948 580224 167000
rect 384672 153144 384724 153196
rect 579620 153144 579672 153196
rect 3240 137844 3292 137896
rect 6276 137844 6328 137896
rect 383108 126896 383160 126948
rect 580172 126896 580224 126948
rect 384580 113092 384632 113144
rect 580172 113092 580224 113144
rect 2780 110712 2832 110764
rect 4988 110712 5040 110764
rect 3332 97860 3384 97912
rect 8024 97860 8076 97912
rect 383016 86912 383068 86964
rect 580172 86912 580224 86964
rect 2780 85008 2832 85060
rect 6184 85008 6236 85060
rect 384396 73108 384448 73160
rect 580172 73108 580224 73160
rect 2780 71612 2832 71664
rect 4896 71612 4948 71664
rect 385684 60664 385736 60716
rect 580172 60664 580224 60716
rect 3056 59304 3108 59356
rect 7840 59304 7892 59356
rect 382924 46860 382976 46912
rect 580172 46860 580224 46912
rect 3424 45500 3476 45552
rect 7748 45500 7800 45552
rect 384488 33056 384540 33108
rect 580172 33056 580224 33108
rect 2780 32988 2832 33040
rect 4804 32988 4856 33040
rect 384304 20612 384356 20664
rect 579988 20612 580040 20664
rect 3056 20136 3108 20188
rect 7656 20136 7708 20188
rect 119896 13472 119948 13524
rect 265164 13472 265216 13524
rect 117228 13404 117280 13456
rect 263784 13404 263836 13456
rect 112812 13336 112864 13388
rect 262496 13336 262548 13388
rect 110328 13268 110380 13320
rect 262588 13268 262640 13320
rect 106188 13200 106240 13252
rect 261024 13200 261076 13252
rect 103428 13132 103480 13184
rect 259736 13132 259788 13184
rect 99288 13064 99340 13116
rect 259644 13064 259696 13116
rect 248420 12520 248472 12572
rect 248696 12520 248748 12572
rect 161296 12384 161348 12436
rect 274916 12384 274968 12436
rect 160100 12316 160152 12368
rect 274824 12316 274876 12368
rect 147588 12248 147640 12300
rect 272156 12248 272208 12300
rect 144828 12180 144880 12232
rect 270868 12180 270920 12232
rect 362500 12180 362552 12232
rect 503720 12180 503772 12232
rect 140044 12112 140096 12164
rect 269488 12112 269540 12164
rect 363972 12112 364024 12164
rect 507216 12112 507268 12164
rect 136456 12044 136508 12096
rect 269396 12044 269448 12096
rect 366732 12044 366784 12096
rect 517888 12044 517940 12096
rect 125876 11976 125928 12028
rect 266636 11976 266688 12028
rect 368112 11976 368164 12028
rect 525432 11976 525484 12028
rect 95148 11908 95200 11960
rect 258356 11908 258408 11960
rect 372344 11908 372396 11960
rect 539600 11908 539652 11960
rect 92388 11840 92440 11892
rect 258264 11840 258316 11892
rect 373540 11840 373592 11892
rect 546684 11840 546736 11892
rect 87972 11772 88024 11824
rect 256976 11772 257028 11824
rect 380532 11772 380584 11824
rect 575112 11772 575164 11824
rect 85488 11704 85540 11756
rect 255412 11704 255464 11756
rect 382004 11704 382056 11756
rect 581000 11704 581052 11756
rect 164884 11636 164936 11688
rect 276388 11636 276440 11688
rect 174268 11568 174320 11620
rect 278964 11568 279016 11620
rect 177856 11500 177908 11552
rect 279056 11500 279108 11552
rect 181444 11432 181496 11484
rect 280528 11432 280580 11484
rect 184940 11364 184992 11416
rect 281816 11364 281868 11416
rect 205548 11296 205600 11348
rect 285956 11296 286008 11348
rect 209044 11228 209096 11280
rect 287428 11228 287480 11280
rect 212172 11160 212224 11212
rect 288716 11160 288768 11212
rect 215668 11092 215720 11144
rect 288624 11092 288676 11144
rect 91008 10956 91060 11008
rect 256884 10956 256936 11008
rect 357072 10956 357124 11008
rect 480536 10956 480588 11008
rect 86684 10888 86736 10940
rect 256792 10888 256844 10940
rect 357348 10888 357400 10940
rect 481640 10888 481692 10940
rect 84108 10820 84160 10872
rect 255596 10820 255648 10872
rect 357256 10820 357308 10872
rect 481732 10820 481784 10872
rect 74448 10752 74500 10804
rect 252744 10752 252796 10804
rect 358728 10752 358780 10804
rect 484768 10752 484820 10804
rect 70308 10684 70360 10736
rect 252836 10684 252888 10736
rect 357164 10684 357216 10736
rect 484032 10684 484084 10736
rect 67548 10616 67600 10668
rect 251456 10616 251508 10668
rect 358452 10616 358504 10668
rect 486424 10616 486476 10668
rect 63224 10548 63276 10600
rect 249892 10548 249944 10600
rect 358544 10548 358596 10600
rect 487160 10548 487212 10600
rect 60648 10480 60700 10532
rect 249984 10480 250036 10532
rect 358636 10480 358688 10532
rect 488816 10480 488868 10532
rect 56508 10412 56560 10464
rect 248420 10412 248472 10464
rect 359924 10412 359976 10464
rect 490012 10412 490064 10464
rect 53656 10344 53708 10396
rect 247316 10344 247368 10396
rect 359740 10344 359792 10396
rect 489920 10344 489972 10396
rect 49608 10276 49660 10328
rect 247408 10276 247460 10328
rect 359832 10276 359884 10328
rect 493048 10276 493100 10328
rect 95056 10208 95108 10260
rect 258172 10208 258224 10260
rect 355784 10208 355836 10260
rect 476488 10208 476540 10260
rect 97908 10140 97960 10192
rect 259552 10140 259604 10192
rect 355692 10140 355744 10192
rect 473452 10140 473504 10192
rect 102048 10072 102100 10124
rect 259828 10072 259880 10124
rect 355876 10072 355928 10124
rect 473360 10072 473412 10124
rect 104532 10004 104584 10056
rect 260932 10004 260984 10056
rect 334992 10004 335044 10056
rect 395344 10004 395396 10056
rect 108948 9936 109000 9988
rect 262312 9936 262364 9988
rect 334900 9936 334952 9988
rect 392584 9936 392636 9988
rect 111616 9868 111668 9920
rect 262404 9868 262456 9920
rect 335084 9868 335136 9920
rect 391112 9868 391164 9920
rect 115848 9800 115900 9852
rect 263692 9800 263744 9852
rect 333704 9800 333756 9852
rect 389456 9800 389508 9852
rect 119804 9732 119856 9784
rect 265256 9732 265308 9784
rect 333612 9732 333664 9784
rect 387800 9732 387852 9784
rect 122748 9664 122800 9716
rect 265072 9664 265124 9716
rect 332140 9664 332192 9716
rect 384304 9664 384356 9716
rect 199108 9596 199160 9648
rect 284576 9596 284628 9648
rect 343272 9596 343324 9648
rect 428464 9596 428516 9648
rect 195612 9528 195664 9580
rect 284668 9528 284720 9580
rect 344652 9528 344704 9580
rect 432052 9528 432104 9580
rect 192024 9460 192076 9512
rect 283288 9460 283340 9512
rect 346032 9460 346084 9512
rect 435548 9460 435600 9512
rect 188528 9392 188580 9444
rect 281724 9392 281776 9444
rect 346124 9392 346176 9444
rect 439136 9392 439188 9444
rect 156604 9324 156656 9376
rect 273628 9324 273680 9376
rect 347412 9324 347464 9376
rect 442632 9324 442684 9376
rect 153016 9256 153068 9308
rect 273536 9256 273588 9308
rect 348884 9256 348936 9308
rect 446220 9256 446272 9308
rect 149520 9188 149572 9240
rect 272064 9188 272116 9240
rect 348976 9188 349028 9240
rect 449808 9188 449860 9240
rect 145932 9120 145984 9172
rect 270776 9120 270828 9172
rect 350264 9120 350316 9172
rect 453304 9120 453356 9172
rect 142436 9052 142488 9104
rect 270684 9052 270736 9104
rect 351552 9052 351604 9104
rect 456892 9052 456944 9104
rect 138848 8984 138900 9036
rect 269212 8984 269264 9036
rect 351644 8984 351696 9036
rect 460388 8984 460440 9036
rect 33600 8916 33652 8968
rect 242992 8916 243044 8968
rect 248788 8916 248840 8968
rect 296904 8916 296956 8968
rect 352840 8916 352892 8968
rect 463976 8916 464028 8968
rect 202696 8848 202748 8900
rect 285864 8848 285916 8900
rect 343364 8848 343416 8900
rect 424968 8848 425020 8900
rect 206192 8780 206244 8832
rect 287244 8780 287296 8832
rect 341984 8780 342036 8832
rect 421380 8780 421432 8832
rect 209780 8712 209832 8764
rect 287336 8712 287388 8764
rect 340604 8712 340656 8764
rect 417884 8712 417936 8764
rect 213368 8644 213420 8696
rect 288532 8644 288584 8696
rect 340696 8644 340748 8696
rect 414296 8644 414348 8696
rect 216864 8576 216916 8628
rect 290004 8576 290056 8628
rect 339132 8576 339184 8628
rect 410800 8576 410852 8628
rect 220452 8508 220504 8560
rect 289912 8508 289964 8560
rect 337752 8508 337804 8560
rect 407212 8508 407264 8560
rect 223948 8440 224000 8492
rect 291568 8440 291620 8492
rect 337844 8440 337896 8492
rect 403532 8440 403584 8492
rect 227536 8372 227588 8424
rect 291476 8372 291528 8424
rect 336372 8372 336424 8424
rect 400128 8372 400180 8424
rect 231032 8304 231084 8356
rect 292856 8304 292908 8356
rect 335176 8304 335228 8356
rect 396540 8304 396592 8356
rect 151820 8236 151872 8288
rect 273352 8236 273404 8288
rect 366824 8236 366876 8288
rect 520740 8236 520792 8288
rect 148324 8168 148376 8220
rect 271972 8168 272024 8220
rect 368204 8168 368256 8220
rect 524236 8168 524288 8220
rect 144736 8100 144788 8152
rect 270592 8100 270644 8152
rect 369492 8100 369544 8152
rect 527824 8100 527876 8152
rect 141240 8032 141292 8084
rect 270500 8032 270552 8084
rect 369584 8032 369636 8084
rect 531320 8032 531372 8084
rect 137652 7964 137704 8016
rect 269120 7964 269172 8016
rect 370872 7964 370924 8016
rect 534908 7964 534960 8016
rect 134156 7896 134208 7948
rect 267924 7896 267976 7948
rect 370964 7896 371016 7948
rect 538404 7896 538456 7948
rect 128176 7828 128228 7880
rect 266544 7828 266596 7880
rect 372436 7828 372488 7880
rect 541992 7828 542044 7880
rect 76196 7760 76248 7812
rect 72608 7692 72660 7744
rect 252652 7760 252704 7812
rect 261760 7760 261812 7812
rect 301044 7760 301096 7812
rect 373632 7760 373684 7812
rect 545488 7760 545540 7812
rect 69112 7624 69164 7676
rect 65524 7556 65576 7608
rect 251364 7692 251416 7744
rect 258264 7692 258316 7744
rect 299572 7692 299624 7744
rect 373724 7692 373776 7744
rect 549076 7692 549128 7744
rect 251272 7624 251324 7676
rect 254676 7624 254728 7676
rect 298284 7624 298336 7676
rect 374920 7624 374972 7676
rect 552664 7624 552716 7676
rect 251180 7556 251232 7608
rect 298376 7556 298428 7608
rect 376484 7556 376536 7608
rect 556160 7556 556212 7608
rect 155408 7488 155460 7540
rect 273444 7488 273496 7540
rect 366916 7488 366968 7540
rect 517152 7488 517204 7540
rect 158904 7420 158956 7472
rect 274732 7420 274784 7472
rect 365444 7420 365496 7472
rect 513564 7420 513616 7472
rect 163688 7352 163740 7404
rect 276296 7352 276348 7404
rect 364064 7352 364116 7404
rect 510068 7352 510120 7404
rect 167184 7284 167236 7336
rect 276204 7284 276256 7336
rect 364156 7284 364208 7336
rect 506480 7284 506532 7336
rect 170772 7216 170824 7268
rect 277584 7216 277636 7268
rect 362684 7216 362736 7268
rect 502984 7216 503036 7268
rect 222752 7148 222804 7200
rect 291384 7148 291436 7200
rect 361396 7148 361448 7200
rect 499396 7148 499448 7200
rect 229836 7080 229888 7132
rect 292764 7080 292816 7132
rect 361304 7080 361356 7132
rect 495900 7080 495952 7132
rect 233424 7012 233476 7064
rect 294328 7012 294380 7064
rect 360108 7012 360160 7064
rect 492312 7012 492364 7064
rect 219256 6944 219308 6996
rect 246304 6944 246356 6996
rect 247592 6944 247644 6996
rect 296812 6944 296864 6996
rect 332232 6944 332284 6996
rect 385960 6944 386012 6996
rect 254032 6876 254084 6928
rect 173164 6808 173216 6860
rect 277676 6808 277728 6860
rect 332324 6808 332376 6860
rect 382372 6808 382424 6860
rect 393964 6808 394016 6860
rect 580172 6808 580224 6860
rect 169576 6740 169628 6792
rect 277492 6740 277544 6792
rect 344744 6740 344796 6792
rect 430856 6740 430908 6792
rect 166080 6672 166132 6724
rect 276112 6672 276164 6724
rect 344836 6672 344888 6724
rect 434444 6672 434496 6724
rect 3424 6604 3476 6656
rect 7564 6604 7616 6656
rect 162492 6604 162544 6656
rect 276020 6604 276072 6656
rect 346216 6604 346268 6656
rect 437940 6604 437992 6656
rect 157800 6536 157852 6588
rect 274640 6536 274692 6588
rect 347504 6536 347556 6588
rect 441528 6536 441580 6588
rect 154212 6468 154264 6520
rect 273260 6468 273312 6520
rect 347596 6468 347648 6520
rect 445024 6468 445076 6520
rect 150624 6400 150676 6452
rect 271880 6400 271932 6452
rect 349068 6400 349120 6452
rect 448612 6400 448664 6452
rect 130568 6332 130620 6384
rect 267832 6332 267884 6384
rect 350448 6332 350500 6384
rect 452108 6332 452160 6384
rect 126980 6264 127032 6316
rect 266452 6264 266504 6316
rect 350356 6264 350408 6316
rect 455696 6264 455748 6316
rect 61936 6196 61988 6248
rect 250076 6196 250128 6248
rect 351736 6196 351788 6248
rect 459192 6196 459244 6248
rect 4068 6128 4120 6180
rect 234896 6128 234948 6180
rect 238116 6128 238168 6180
rect 294236 6128 294288 6180
rect 353116 6128 353168 6180
rect 462780 6128 462832 6180
rect 176660 6060 176712 6112
rect 278872 6060 278924 6112
rect 343456 6060 343508 6112
rect 427268 6060 427320 6112
rect 180248 5992 180300 6044
rect 280344 5992 280396 6044
rect 342076 5992 342128 6044
rect 423772 5992 423824 6044
rect 183744 5924 183796 5976
rect 280436 5924 280488 5976
rect 342168 5924 342220 5976
rect 420184 5924 420236 5976
rect 187332 5856 187384 5908
rect 281632 5856 281684 5908
rect 340788 5856 340840 5908
rect 416688 5856 416740 5908
rect 190828 5788 190880 5840
rect 283196 5788 283248 5840
rect 339316 5788 339368 5840
rect 413100 5788 413152 5840
rect 194416 5720 194468 5772
rect 283104 5720 283156 5772
rect 339224 5720 339276 5772
rect 409604 5720 409656 5772
rect 197912 5652 197964 5704
rect 284484 5652 284536 5704
rect 338028 5652 338080 5704
rect 406016 5652 406068 5704
rect 201500 5584 201552 5636
rect 285772 5584 285824 5636
rect 337936 5584 337988 5636
rect 402520 5584 402572 5636
rect 226340 5516 226392 5568
rect 291292 5516 291344 5568
rect 336464 5516 336516 5568
rect 398932 5516 398984 5568
rect 203892 5448 203944 5500
rect 285680 5448 285732 5500
rect 326712 5448 326764 5500
rect 359924 5448 359976 5500
rect 368388 5448 368440 5500
rect 526628 5448 526680 5500
rect 200304 5380 200356 5432
rect 284392 5380 284444 5432
rect 326804 5380 326856 5432
rect 361120 5380 361172 5432
rect 369676 5380 369728 5432
rect 530124 5380 530176 5432
rect 123484 5312 123536 5364
rect 191104 5312 191156 5364
rect 193220 5312 193272 5364
rect 124680 5244 124732 5296
rect 193864 5244 193916 5296
rect 196808 5312 196860 5364
rect 284300 5312 284352 5364
rect 328092 5312 328144 5364
rect 364616 5312 364668 5364
rect 371056 5312 371108 5364
rect 533712 5312 533764 5364
rect 283012 5244 283064 5296
rect 326620 5244 326672 5296
rect 363512 5244 363564 5296
rect 371148 5244 371200 5296
rect 537208 5244 537260 5296
rect 189724 5176 189776 5228
rect 282920 5176 282972 5228
rect 328000 5176 328052 5228
rect 367008 5176 367060 5228
rect 372528 5176 372580 5228
rect 540796 5176 540848 5228
rect 186136 5108 186188 5160
rect 281540 5108 281592 5160
rect 328184 5108 328236 5160
rect 368204 5108 368256 5160
rect 373908 5108 373960 5160
rect 544384 5108 544436 5160
rect 182548 5040 182600 5092
rect 280252 5040 280304 5092
rect 329656 5040 329708 5092
rect 370596 5040 370648 5092
rect 373816 5040 373868 5092
rect 547880 5040 547932 5092
rect 179052 4972 179104 5024
rect 280160 4972 280212 5024
rect 329472 4972 329524 5024
rect 371700 4972 371752 5024
rect 375012 4972 375064 5024
rect 551468 4972 551520 5024
rect 7656 4904 7708 4956
rect 234620 4904 234672 4956
rect 2872 4836 2924 4888
rect 234712 4836 234764 4888
rect 236092 4836 236144 4888
rect 237012 4836 237064 4888
rect 271236 4904 271288 4956
rect 302424 4904 302476 4956
rect 329564 4904 329616 4956
rect 374092 4904 374144 4956
rect 375104 4904 375156 4956
rect 554964 4904 555016 4956
rect 294052 4836 294104 4888
rect 330852 4836 330904 4888
rect 377680 4836 377732 4888
rect 378048 4836 378100 4888
rect 562048 4836 562100 4888
rect 1676 4768 1728 4820
rect 232228 4768 232280 4820
rect 244924 4768 244976 4820
rect 294144 4768 294196 4820
rect 330760 4768 330812 4820
rect 378876 4768 378928 4820
rect 379336 4768 379388 4820
rect 569132 4768 569184 4820
rect 207388 4700 207440 4752
rect 287060 4700 287112 4752
rect 325424 4700 325476 4752
rect 357532 4700 357584 4752
rect 368296 4700 368348 4752
rect 523040 4700 523092 4752
rect 210976 4632 211028 4684
rect 287152 4632 287204 4684
rect 325516 4632 325568 4684
rect 356336 4632 356388 4684
rect 366916 4632 366968 4684
rect 519544 4632 519596 4684
rect 214472 4564 214524 4616
rect 288440 4564 288492 4616
rect 325332 4564 325384 4616
rect 354036 4564 354088 4616
rect 365628 4564 365680 4616
rect 515956 4564 516008 4616
rect 171968 4496 172020 4548
rect 245016 4496 245068 4548
rect 274824 4496 274876 4548
rect 303804 4496 303856 4548
rect 323952 4496 324004 4548
rect 352840 4496 352892 4548
rect 365536 4496 365588 4548
rect 512460 4496 512512 4548
rect 221556 4428 221608 4480
rect 290096 4428 290148 4480
rect 323860 4428 323912 4480
rect 349252 4428 349304 4480
rect 364248 4428 364300 4480
rect 508872 4428 508924 4480
rect 225144 4360 225196 4412
rect 291200 4360 291252 4412
rect 322664 4360 322716 4412
rect 345756 4360 345808 4412
rect 362776 4360 362828 4412
rect 505376 4360 505428 4412
rect 228732 4292 228784 4344
rect 292672 4292 292724 4344
rect 362868 4292 362920 4344
rect 501788 4292 501840 4344
rect 234804 4224 234856 4276
rect 235816 4224 235868 4276
rect 143540 4156 143592 4208
rect 144828 4156 144880 4208
rect 218060 4156 218112 4208
rect 292580 4224 292632 4276
rect 361488 4224 361540 4276
rect 498200 4224 498252 4276
rect 293960 4156 294012 4208
rect 332416 4156 332468 4208
rect 381176 4156 381228 4208
rect 489920 4156 489972 4208
rect 491116 4156 491168 4208
rect 50160 4088 50212 4140
rect 46664 4020 46716 4072
rect 245936 4088 245988 4140
rect 279516 4088 279568 4140
rect 305276 4088 305328 4140
rect 307944 4088 307996 4140
rect 328368 4088 328420 4140
rect 332508 4088 332560 4140
rect 244096 4020 244148 4072
rect 249064 4020 249116 4072
rect 276020 4020 276072 4072
rect 303896 4020 303948 4072
rect 320088 4020 320140 4072
rect 333888 4020 333940 4072
rect 365812 4088 365864 4140
rect 396724 4088 396776 4140
rect 521844 4088 521896 4140
rect 45376 3952 45428 4004
rect 245752 3952 245804 4004
rect 277124 3952 277176 4004
rect 305092 3952 305144 4004
rect 324964 3952 325016 4004
rect 332692 3952 332744 4004
rect 39580 3884 39632 3936
rect 244372 3884 244424 3936
rect 265348 3884 265400 3936
rect 271144 3884 271196 3936
rect 272432 3884 272484 3936
rect 303712 3884 303764 3936
rect 305552 3884 305604 3936
rect 311992 3884 312044 3936
rect 326988 3884 327040 3936
rect 331128 3884 331180 3936
rect 376484 4020 376536 4072
rect 399484 4020 399536 4072
rect 529020 4020 529072 4072
rect 379980 3952 380032 4004
rect 405004 3952 405056 4004
rect 536104 3952 536156 4004
rect 383568 3884 383620 3936
rect 403624 3884 403676 3936
rect 543188 3884 543240 3936
rect 35992 3816 36044 3868
rect 37096 3816 37148 3868
rect 38384 3816 38436 3868
rect 244648 3816 244700 3868
rect 270040 3816 270092 3868
rect 302332 3816 302384 3868
rect 304356 3816 304408 3868
rect 311164 3816 311216 3868
rect 320824 3816 320876 3868
rect 326804 3816 326856 3868
rect 328276 3816 328328 3868
rect 333796 3816 333848 3868
rect 387156 3816 387208 3868
rect 411904 3816 411956 3868
rect 557356 3816 557408 3868
rect 31300 3748 31352 3800
rect 241888 3748 241940 3800
rect 264152 3748 264204 3800
rect 301136 3748 301188 3800
rect 301964 3748 302016 3800
rect 310796 3748 310848 3800
rect 322204 3748 322256 3800
rect 330392 3748 330444 3800
rect 32404 3680 32456 3732
rect 243084 3680 243136 3732
rect 245200 3680 245252 3732
rect 254584 3680 254636 3732
rect 257068 3680 257120 3732
rect 299664 3680 299716 3732
rect 305460 3680 305512 3732
rect 310704 3680 310756 3732
rect 321284 3680 321336 3732
rect 342168 3748 342220 3800
rect 343548 3748 343600 3800
rect 426164 3748 426216 3800
rect 333704 3680 333756 3732
rect 390652 3680 390704 3732
rect 391204 3680 391256 3732
rect 415492 3680 415544 3732
rect 416044 3680 416096 3732
rect 422576 3680 422628 3732
rect 425704 3680 425756 3732
rect 429844 3748 429896 3800
rect 432512 3748 432564 3800
rect 432604 3748 432656 3800
rect 440332 3748 440384 3800
rect 571524 3748 571576 3800
rect 564440 3680 564492 3732
rect 28816 3612 28868 3664
rect 241612 3612 241664 3664
rect 241704 3612 241756 3664
rect 251824 3612 251876 3664
rect 253480 3612 253532 3664
rect 298468 3612 298520 3664
rect 298560 3612 298612 3664
rect 309140 3612 309192 3664
rect 321376 3612 321428 3664
rect 337476 3612 337528 3664
rect 338764 3612 338816 3664
rect 404820 3612 404872 3664
rect 413284 3612 413336 3664
rect 560852 3612 560904 3664
rect 11152 3544 11204 3596
rect 12348 3544 12400 3596
rect 25320 3544 25372 3596
rect 240508 3544 240560 3596
rect 247040 3544 247092 3596
rect 255872 3544 255924 3596
rect 256608 3544 256660 3596
rect 298192 3544 298244 3596
rect 300768 3544 300820 3596
rect 572 3476 624 3528
rect 1308 3476 1360 3528
rect 9956 3476 10008 3528
rect 10968 3476 11020 3528
rect 18236 3476 18288 3528
rect 19248 3476 19300 3528
rect 24216 3476 24268 3528
rect 240324 3476 240376 3528
rect 246396 3476 246448 3528
rect 296996 3476 297048 3528
rect 297272 3476 297324 3528
rect 309324 3544 309376 3596
rect 317328 3544 317380 3596
rect 325516 3544 325568 3596
rect 327724 3544 327776 3596
rect 331588 3544 331640 3596
rect 369400 3544 369452 3596
rect 369768 3544 369820 3596
rect 532516 3544 532568 3596
rect 306748 3476 306800 3528
rect 307668 3476 307720 3528
rect 23020 3408 23072 3460
rect 240232 3408 240284 3460
rect 242900 3408 242952 3460
rect 27712 3340 27764 3392
rect 28908 3340 28960 3392
rect 34796 3340 34848 3392
rect 35808 3340 35860 3392
rect 40684 3340 40736 3392
rect 41328 3340 41380 3392
rect 41880 3340 41932 3392
rect 42708 3340 42760 3392
rect 43076 3340 43128 3392
rect 44088 3340 44140 3392
rect 44272 3340 44324 3392
rect 45468 3340 45520 3392
rect 48964 3340 49016 3392
rect 49608 3340 49660 3392
rect 52552 3340 52604 3392
rect 53656 3340 53708 3392
rect 56048 3340 56100 3392
rect 56508 3340 56560 3392
rect 59636 3340 59688 3392
rect 60648 3340 60700 3392
rect 60832 3340 60884 3392
rect 62028 3340 62080 3392
rect 66720 3340 66772 3392
rect 67548 3340 67600 3392
rect 67916 3340 67968 3392
rect 68928 3340 68980 3392
rect 57244 3272 57296 3324
rect 248696 3340 248748 3392
rect 249984 3340 250036 3392
rect 259460 3340 259512 3392
rect 260748 3340 260800 3392
rect 273628 3340 273680 3392
rect 274548 3340 274600 3392
rect 278320 3408 278372 3460
rect 282184 3408 282236 3460
rect 284300 3408 284352 3460
rect 285588 3408 285640 3460
rect 287796 3408 287848 3460
rect 288348 3408 288400 3460
rect 288992 3408 289044 3460
rect 289728 3408 289780 3460
rect 295708 3408 295760 3460
rect 296076 3408 296128 3460
rect 309232 3476 309284 3528
rect 313280 3476 313332 3528
rect 313832 3476 313884 3528
rect 320916 3476 320968 3528
rect 322112 3476 322164 3528
rect 322296 3476 322348 3528
rect 323308 3476 323360 3528
rect 309048 3408 309100 3460
rect 312176 3408 312228 3460
rect 299664 3340 299716 3392
rect 64328 3204 64380 3256
rect 251548 3272 251600 3324
rect 283104 3272 283156 3324
rect 73804 3204 73856 3256
rect 74448 3204 74500 3256
rect 75000 3204 75052 3256
rect 75828 3204 75880 3256
rect 77392 3204 77444 3256
rect 78588 3204 78640 3256
rect 80888 3204 80940 3256
rect 81348 3204 81400 3256
rect 82084 3204 82136 3256
rect 82728 3204 82780 3256
rect 84476 3204 84528 3256
rect 85488 3204 85540 3256
rect 85672 3204 85724 3256
rect 86776 3204 86828 3256
rect 90364 3204 90416 3256
rect 91008 3204 91060 3256
rect 91560 3204 91612 3256
rect 92388 3204 92440 3256
rect 71504 3136 71556 3188
rect 252928 3204 252980 3256
rect 281908 3204 281960 3256
rect 307944 3340 307996 3392
rect 312084 3340 312136 3392
rect 318616 3340 318668 3392
rect 328000 3476 328052 3528
rect 331036 3476 331088 3528
rect 372896 3476 372948 3528
rect 375196 3476 375248 3528
rect 550272 3476 550324 3528
rect 329196 3408 329248 3460
rect 330944 3408 330996 3460
rect 375288 3408 375340 3460
rect 375380 3408 375432 3460
rect 553768 3408 553820 3460
rect 324228 3340 324280 3392
rect 351644 3340 351696 3392
rect 354588 3340 354640 3392
rect 472256 3340 472308 3392
rect 473360 3340 473412 3392
rect 474556 3340 474608 3392
rect 481640 3340 481692 3392
rect 482836 3340 482888 3392
rect 310612 3272 310664 3324
rect 311440 3272 311492 3324
rect 313372 3272 313424 3324
rect 318708 3272 318760 3324
rect 329748 3272 329800 3324
rect 362316 3272 362368 3324
rect 398104 3272 398156 3324
rect 514760 3272 514812 3324
rect 83280 3068 83332 3120
rect 84108 3068 84160 3120
rect 78588 3000 78640 3052
rect 254308 3136 254360 3188
rect 266544 3136 266596 3188
rect 267648 3136 267700 3188
rect 285404 3136 285456 3188
rect 92756 3068 92808 3120
rect 93768 3068 93820 3120
rect 93952 3068 94004 3120
rect 95056 3068 95108 3120
rect 97448 3068 97500 3120
rect 97908 3068 97960 3120
rect 98644 3068 98696 3120
rect 99288 3068 99340 3120
rect 99840 3068 99892 3120
rect 100668 3068 100720 3120
rect 256700 3068 256752 3120
rect 280712 3068 280764 3120
rect 89168 2932 89220 2984
rect 96252 2932 96304 2984
rect 258448 3000 258500 3052
rect 290188 3000 290240 3052
rect 305184 3136 305236 3188
rect 324044 3204 324096 3256
rect 350448 3204 350500 3256
rect 353208 3204 353260 3256
rect 465172 3204 465224 3256
rect 306472 3136 306524 3188
rect 324136 3136 324188 3188
rect 348056 3136 348108 3188
rect 351828 3136 351880 3188
rect 458088 3136 458140 3188
rect 306564 3068 306616 3120
rect 318156 3068 318208 3120
rect 320916 3068 320968 3120
rect 322848 3068 322900 3120
rect 344560 3068 344612 3120
rect 347688 3068 347740 3120
rect 443828 3068 443880 3120
rect 443920 3068 443972 3120
rect 293684 3000 293736 3052
rect 309416 3000 309468 3052
rect 310244 3000 310296 3052
rect 313464 3000 313516 3052
rect 322756 3000 322808 3052
rect 343364 3000 343416 3052
rect 346308 3000 346360 3052
rect 436744 3000 436796 3052
rect 440884 3000 440936 3052
rect 454500 3068 454552 3120
rect 102232 2932 102284 2984
rect 103428 2932 103480 2984
rect 105728 2932 105780 2984
rect 106188 2932 106240 2984
rect 106924 2932 106976 2984
rect 107568 2932 107620 2984
rect 108120 2932 108172 2984
rect 108948 2932 109000 2984
rect 109316 2932 109368 2984
rect 110328 2932 110380 2984
rect 101036 2864 101088 2916
rect 102048 2864 102100 2916
rect 103336 2864 103388 2916
rect 261116 2932 261168 2984
rect 291384 2932 291436 2984
rect 307852 2932 307904 2984
rect 321468 2932 321520 2984
rect 340972 2932 341024 2984
rect 344928 2932 344980 2984
rect 429660 2932 429712 2984
rect 110512 2864 110564 2916
rect 262680 2864 262732 2916
rect 262956 2864 263008 2916
rect 263508 2864 263560 2916
rect 294880 2864 294932 2916
rect 309508 2864 309560 2916
rect 312636 2864 312688 2916
rect 313556 2864 313608 2916
rect 317236 2864 317288 2916
rect 324412 2864 324464 2916
rect 326896 2864 326948 2916
rect 114008 2796 114060 2848
rect 114468 2796 114520 2848
rect 115204 2796 115256 2848
rect 115848 2796 115900 2848
rect 116400 2796 116452 2848
rect 117228 2796 117280 2848
rect 117596 2796 117648 2848
rect 118792 2796 118844 2848
rect 119804 2796 119856 2848
rect 263876 2796 263928 2848
rect 292580 2796 292632 2848
rect 308220 2796 308272 2848
rect 325608 2796 325660 2848
rect 358728 2864 358780 2916
rect 383200 2864 383252 2916
rect 408408 2864 408460 2916
rect 417424 2864 417476 2916
rect 355232 2796 355284 2848
rect 405096 2796 405148 2848
rect 418620 2796 418672 2848
rect 418804 2864 418856 2916
rect 425796 2728 425848 2780
rect 432512 2864 432564 2916
rect 433248 2864 433300 2916
rect 436928 2932 436980 2984
rect 447416 2932 447468 2984
rect 447784 3000 447836 3052
rect 468668 3000 468720 3052
rect 461584 2932 461636 2984
rect 479340 2864 479392 2916
rect 450912 2796 450964 2848
rect 451004 2796 451056 2848
rect 475752 2796 475804 2848
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 284036 703582 284248 703610
rect 8128 700369 8156 703520
rect 24320 700505 24348 703520
rect 40512 700641 40540 703520
rect 40498 700632 40554 700641
rect 40498 700567 40554 700576
rect 24306 700496 24362 700505
rect 24306 700431 24362 700440
rect 8114 700360 8170 700369
rect 72988 700330 73016 703520
rect 89180 700534 89208 703520
rect 105464 700602 105492 703520
rect 137848 700738 137876 703520
rect 154132 700942 154160 703520
rect 170324 701010 170352 703520
rect 170312 701004 170364 701010
rect 170312 700946 170364 700952
rect 154120 700936 154172 700942
rect 154120 700878 154172 700884
rect 137836 700732 137888 700738
rect 137836 700674 137888 700680
rect 105452 700596 105504 700602
rect 105452 700538 105504 700544
rect 89168 700528 89220 700534
rect 89168 700470 89220 700476
rect 8114 700295 8170 700304
rect 72976 700324 73028 700330
rect 72976 700266 73028 700272
rect 202800 700194 202828 703520
rect 218992 702434 219020 703520
rect 218992 702406 219388 702434
rect 202788 700188 202840 700194
rect 202788 700130 202840 700136
rect 3422 684312 3478 684321
rect 3422 684247 3478 684256
rect 3436 683194 3464 684247
rect 3424 683188 3476 683194
rect 3424 683130 3476 683136
rect 3514 671256 3570 671265
rect 3514 671191 3570 671200
rect 3528 670750 3556 671191
rect 3516 670744 3568 670750
rect 3516 670686 3568 670692
rect 3422 658200 3478 658209
rect 3422 658135 3478 658144
rect 3436 656946 3464 658135
rect 3424 656940 3476 656946
rect 3424 656882 3476 656888
rect 3424 632120 3476 632126
rect 3422 632088 3424 632097
rect 3476 632088 3478 632097
rect 3422 632023 3478 632032
rect 3146 619168 3202 619177
rect 3146 619103 3202 619112
rect 3160 618322 3188 619103
rect 3148 618316 3200 618322
rect 3148 618258 3200 618264
rect 3238 606112 3294 606121
rect 3238 606047 3294 606056
rect 3252 605878 3280 606047
rect 3240 605872 3292 605878
rect 3240 605814 3292 605820
rect 3330 580000 3386 580009
rect 3330 579935 3386 579944
rect 3344 579698 3372 579935
rect 3332 579692 3384 579698
rect 3332 579634 3384 579640
rect 3422 566944 3478 566953
rect 3422 566879 3478 566888
rect 3436 565894 3464 566879
rect 3424 565888 3476 565894
rect 3424 565830 3476 565836
rect 3422 553888 3478 553897
rect 3422 553823 3478 553832
rect 3436 553450 3464 553823
rect 3424 553444 3476 553450
rect 3424 553386 3476 553392
rect 3422 527912 3478 527921
rect 3422 527847 3478 527856
rect 3436 527202 3464 527847
rect 3424 527196 3476 527202
rect 3424 527138 3476 527144
rect 3422 514856 3478 514865
rect 3422 514791 3424 514800
rect 3476 514791 3478 514800
rect 3424 514762 3476 514768
rect 3054 501800 3110 501809
rect 3054 501735 3110 501744
rect 3068 501022 3096 501735
rect 3056 501016 3108 501022
rect 3056 500958 3108 500964
rect 219360 491094 219388 702406
rect 235184 699990 235212 703520
rect 235172 699984 235224 699990
rect 235172 699926 235224 699932
rect 267660 699854 267688 703520
rect 283852 703474 283880 703520
rect 284036 703474 284064 703582
rect 283852 703446 284064 703474
rect 267648 699848 267700 699854
rect 267648 699790 267700 699796
rect 284116 590708 284168 590714
rect 284116 590650 284168 590656
rect 282828 563100 282880 563106
rect 282828 563042 282880 563048
rect 280068 536852 280120 536858
rect 280068 536794 280120 536800
rect 278688 510672 278740 510678
rect 278688 510614 278740 510620
rect 219348 491088 219400 491094
rect 219348 491030 219400 491036
rect 273168 491020 273220 491026
rect 273168 490962 273220 490968
rect 271788 490952 271840 490958
rect 271788 490894 271840 490900
rect 7932 490884 7984 490890
rect 7932 490826 7984 490832
rect 5448 490816 5500 490822
rect 5448 490758 5500 490764
rect 5356 490748 5408 490754
rect 5356 490690 5408 490696
rect 5264 490680 5316 490686
rect 5264 490622 5316 490628
rect 3332 490612 3384 490618
rect 3332 490554 3384 490560
rect 2780 475720 2832 475726
rect 2778 475688 2780 475697
rect 2832 475688 2834 475697
rect 2778 475623 2834 475632
rect 3240 462732 3292 462738
rect 3240 462674 3292 462680
rect 3252 462641 3280 462674
rect 3238 462632 3294 462641
rect 3238 462567 3294 462576
rect 3240 449608 3292 449614
rect 3238 449576 3240 449585
rect 3292 449576 3294 449585
rect 3238 449511 3294 449520
rect 2780 423632 2832 423638
rect 2778 423600 2780 423609
rect 2832 423600 2834 423609
rect 2778 423535 2834 423544
rect 3344 410553 3372 490554
rect 4068 490544 4120 490550
rect 4068 490486 4120 490492
rect 3976 490476 4028 490482
rect 3976 490418 4028 490424
rect 3884 490340 3936 490346
rect 3884 490282 3936 490288
rect 3792 490204 3844 490210
rect 3792 490146 3844 490152
rect 3608 490068 3660 490074
rect 3608 490010 3660 490016
rect 3424 489932 3476 489938
rect 3424 489874 3476 489880
rect 3330 410544 3386 410553
rect 3330 410479 3386 410488
rect 2780 397588 2832 397594
rect 2780 397530 2832 397536
rect 2792 397497 2820 397530
rect 2778 397488 2834 397497
rect 2778 397423 2834 397432
rect 2780 371476 2832 371482
rect 2780 371418 2832 371424
rect 2792 371385 2820 371418
rect 2778 371376 2834 371385
rect 2778 371311 2834 371320
rect 2780 319864 2832 319870
rect 2780 319806 2832 319812
rect 2792 319297 2820 319806
rect 2778 319288 2834 319297
rect 2778 319223 2834 319232
rect 3148 293820 3200 293826
rect 3148 293762 3200 293768
rect 3160 293185 3188 293762
rect 3146 293176 3202 293185
rect 3146 293111 3202 293120
rect 2780 267300 2832 267306
rect 2780 267242 2832 267248
rect 2792 267209 2820 267242
rect 2778 267200 2834 267209
rect 2778 267135 2834 267144
rect 3240 241120 3292 241126
rect 3238 241088 3240 241097
rect 3292 241088 3294 241097
rect 3238 241023 3294 241032
rect 3240 188896 3292 188902
rect 3238 188864 3240 188873
rect 3292 188864 3294 188873
rect 3238 188799 3294 188808
rect 3436 149841 3464 489874
rect 3516 485852 3568 485858
rect 3516 485794 3568 485800
rect 3528 162897 3556 485794
rect 3620 201929 3648 490010
rect 3700 485920 3752 485926
rect 3700 485862 3752 485868
rect 3712 214985 3740 485862
rect 3804 254153 3832 490146
rect 3896 306241 3924 490282
rect 3988 345409 4016 490418
rect 4080 358465 4108 490486
rect 4712 487620 4764 487626
rect 4712 487562 4764 487568
rect 4724 475726 4752 487562
rect 4988 487552 5040 487558
rect 4988 487494 5040 487500
rect 4896 487416 4948 487422
rect 4896 487358 4948 487364
rect 4804 487212 4856 487218
rect 4804 487154 4856 487160
rect 4712 475720 4764 475726
rect 4712 475662 4764 475668
rect 4066 358456 4122 358465
rect 4066 358391 4122 358400
rect 3974 345400 4030 345409
rect 3974 345335 4030 345344
rect 3882 306232 3938 306241
rect 3882 306167 3938 306176
rect 3790 254144 3846 254153
rect 3790 254079 3846 254088
rect 3698 214976 3754 214985
rect 3698 214911 3754 214920
rect 3606 201920 3662 201929
rect 3606 201855 3662 201864
rect 3514 162888 3570 162897
rect 3514 162823 3570 162832
rect 3422 149832 3478 149841
rect 3422 149767 3478 149776
rect 3240 137896 3292 137902
rect 3240 137838 3292 137844
rect 3252 136785 3280 137838
rect 3238 136776 3294 136785
rect 3238 136711 3294 136720
rect 2780 110764 2832 110770
rect 2780 110706 2832 110712
rect 2792 110673 2820 110706
rect 2778 110664 2834 110673
rect 2778 110599 2834 110608
rect 3332 97912 3384 97918
rect 3332 97854 3384 97860
rect 3344 97617 3372 97854
rect 3330 97608 3386 97617
rect 3330 97543 3386 97552
rect 2780 85060 2832 85066
rect 2780 85002 2832 85008
rect 2792 84697 2820 85002
rect 2778 84688 2834 84697
rect 2778 84623 2834 84632
rect 2780 71664 2832 71670
rect 2778 71632 2780 71641
rect 2832 71632 2834 71641
rect 2778 71567 2834 71576
rect 3056 59356 3108 59362
rect 3056 59298 3108 59304
rect 3068 58585 3096 59298
rect 3054 58576 3110 58585
rect 3054 58511 3110 58520
rect 3424 45552 3476 45558
rect 3422 45520 3424 45529
rect 3476 45520 3478 45529
rect 3422 45455 3478 45464
rect 4816 33046 4844 487154
rect 4908 71670 4936 487358
rect 5000 110770 5028 487494
rect 5172 486056 5224 486062
rect 5172 485998 5224 486004
rect 5080 485988 5132 485994
rect 5080 485930 5132 485936
rect 5092 267306 5120 485930
rect 5184 319870 5212 485998
rect 5276 371482 5304 490622
rect 5368 397594 5396 490690
rect 5460 423638 5488 490758
rect 6552 490408 6604 490414
rect 6552 490350 6604 490356
rect 6460 490272 6512 490278
rect 6460 490214 6512 490220
rect 6368 490136 6420 490142
rect 6368 490078 6420 490084
rect 6276 490000 6328 490006
rect 6276 489942 6328 489948
rect 6182 486024 6238 486033
rect 6182 485959 6238 485968
rect 5448 423632 5500 423638
rect 5448 423574 5500 423580
rect 5356 397588 5408 397594
rect 5356 397530 5408 397536
rect 5264 371476 5316 371482
rect 5264 371418 5316 371424
rect 5446 336016 5502 336025
rect 5446 335951 5502 335960
rect 5172 319864 5224 319870
rect 5172 319806 5224 319812
rect 5080 267300 5132 267306
rect 5080 267242 5132 267248
rect 4988 110764 5040 110770
rect 4988 110706 5040 110712
rect 4896 71664 4948 71670
rect 4896 71606 4948 71612
rect 2780 33040 2832 33046
rect 2780 32982 2832 32988
rect 4804 33040 4856 33046
rect 4804 32982 4856 32988
rect 2792 32473 2820 32982
rect 2778 32464 2834 32473
rect 2778 32399 2834 32408
rect 3056 20188 3108 20194
rect 3056 20130 3108 20136
rect 3068 19417 3096 20130
rect 3054 19408 3110 19417
rect 3054 19343 3110 19352
rect 1306 11656 1362 11665
rect 1306 11591 1362 11600
rect 1320 3534 1348 11591
rect 5460 6914 5488 335951
rect 6196 85066 6224 485959
rect 6288 137902 6316 489942
rect 6380 188902 6408 490078
rect 6472 241126 6500 490214
rect 6564 293826 6592 490350
rect 7748 487484 7800 487490
rect 7748 487426 7800 487432
rect 7564 487348 7616 487354
rect 7564 487290 7616 487296
rect 6644 486124 6696 486130
rect 6644 486066 6696 486072
rect 6656 449614 6684 486066
rect 6644 449608 6696 449614
rect 6644 449550 6696 449556
rect 6552 293820 6604 293826
rect 6552 293762 6604 293768
rect 6460 241120 6512 241126
rect 6460 241062 6512 241068
rect 6368 188896 6420 188902
rect 6368 188838 6420 188844
rect 6276 137896 6328 137902
rect 6276 137838 6328 137844
rect 6184 85060 6236 85066
rect 6184 85002 6236 85008
rect 5276 6886 5488 6914
rect 3424 6656 3476 6662
rect 3424 6598 3476 6604
rect 3436 6497 3464 6598
rect 3422 6488 3478 6497
rect 3422 6423 3478 6432
rect 4068 6180 4120 6186
rect 4068 6122 4120 6128
rect 2872 4888 2924 4894
rect 2872 4830 2924 4836
rect 1676 4820 1728 4826
rect 1676 4762 1728 4768
rect 572 3528 624 3534
rect 572 3470 624 3476
rect 1308 3528 1360 3534
rect 1308 3470 1360 3476
rect 584 480 612 3470
rect 1688 480 1716 4762
rect 2884 480 2912 4830
rect 4080 480 4108 6122
rect 5276 480 5304 6886
rect 7576 6662 7604 487290
rect 7656 487280 7708 487286
rect 7656 487222 7708 487228
rect 7668 20194 7696 487222
rect 7760 45558 7788 487426
rect 7838 485888 7894 485897
rect 7838 485823 7894 485832
rect 7852 59362 7880 485823
rect 7944 462738 7972 490826
rect 242438 490240 242494 490249
rect 242438 490175 242494 490184
rect 238574 490104 238630 490113
rect 238574 490039 238630 490048
rect 237286 489968 237342 489977
rect 237286 489903 237342 489912
rect 235908 487824 235960 487830
rect 235908 487766 235960 487772
rect 235920 487506 235948 487766
rect 237300 487506 237328 489903
rect 238588 487506 238616 490039
rect 239864 487892 239916 487898
rect 239864 487834 239916 487840
rect 239876 487506 239904 487834
rect 242452 487506 242480 490175
rect 268292 488300 268344 488306
rect 268292 488242 268344 488248
rect 255228 488232 255280 488238
rect 255228 488174 255280 488180
rect 247592 488164 247644 488170
rect 247592 488106 247644 488112
rect 243728 488028 243780 488034
rect 243728 487970 243780 487976
rect 243740 487506 243768 487970
rect 245016 487960 245068 487966
rect 245016 487902 245068 487908
rect 245028 487506 245056 487902
rect 247604 487506 247632 488106
rect 248880 488096 248932 488102
rect 248880 488038 248932 488044
rect 248892 487506 248920 488038
rect 250168 487688 250220 487694
rect 250168 487630 250220 487636
rect 250180 487506 250208 487630
rect 255240 487506 255268 488174
rect 268304 487506 268332 488242
rect 269258 487756 269310 487762
rect 269258 487698 269310 487704
rect 235704 487478 235948 487506
rect 236992 487478 237328 487506
rect 238280 487478 238616 487506
rect 239568 487478 239904 487506
rect 242144 487478 242480 487506
rect 243432 487478 243768 487506
rect 244720 487478 245056 487506
rect 247296 487478 247632 487506
rect 248584 487478 248920 487506
rect 249872 487478 250208 487506
rect 255024 487478 255268 487506
rect 267996 487478 268332 487506
rect 269270 487492 269298 487698
rect 271800 487506 271828 490894
rect 273180 487778 273208 490962
rect 275928 488504 275980 488510
rect 275928 488446 275980 488452
rect 274548 488436 274600 488442
rect 274548 488378 274600 488384
rect 273134 487750 273208 487778
rect 271800 487478 271860 487506
rect 273134 487492 273162 487750
rect 274560 487506 274588 488378
rect 275940 487506 275968 488446
rect 277124 488368 277176 488374
rect 277124 488310 277176 488316
rect 277136 487506 277164 488310
rect 278700 487506 278728 510614
rect 280080 487506 280108 536794
rect 281448 524476 281500 524482
rect 281448 524418 281500 524424
rect 281460 489914 281488 524418
rect 282840 489914 282868 563042
rect 284128 489914 284156 590650
rect 284220 491230 284248 703582
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 299388 700868 299440 700874
rect 299388 700810 299440 700816
rect 293866 700768 293922 700777
rect 293866 700703 293922 700712
rect 292488 696992 292540 696998
rect 292488 696934 292540 696940
rect 292396 683256 292448 683262
rect 292396 683198 292448 683204
rect 291108 670812 291160 670818
rect 291108 670754 291160 670760
rect 288348 643136 288400 643142
rect 288348 643078 288400 643084
rect 286968 616888 287020 616894
rect 286968 616830 287020 616836
rect 285588 576904 285640 576910
rect 285588 576846 285640 576852
rect 285600 491298 285628 576846
rect 286980 491298 287008 616830
rect 288360 491298 288388 643078
rect 289728 630692 289780 630698
rect 289728 630634 289780 630640
rect 289740 491298 289768 630634
rect 291120 491298 291148 670754
rect 285128 491292 285180 491298
rect 285128 491234 285180 491240
rect 285588 491292 285640 491298
rect 285588 491234 285640 491240
rect 286416 491292 286468 491298
rect 286416 491234 286468 491240
rect 286968 491292 287020 491298
rect 286968 491234 287020 491240
rect 287704 491292 287756 491298
rect 287704 491234 287756 491240
rect 288348 491292 288400 491298
rect 288348 491234 288400 491240
rect 288992 491292 289044 491298
rect 288992 491234 289044 491240
rect 289728 491292 289780 491298
rect 289728 491234 289780 491240
rect 290280 491292 290332 491298
rect 290280 491234 290332 491240
rect 291108 491292 291160 491298
rect 291108 491234 291160 491240
rect 291568 491292 291620 491298
rect 291568 491234 291620 491240
rect 284208 491224 284260 491230
rect 284208 491166 284260 491172
rect 281368 489886 281488 489914
rect 282656 489886 282868 489914
rect 283944 489886 284156 489914
rect 281368 487506 281396 489886
rect 282656 487506 282684 489886
rect 283944 487506 283972 489886
rect 285140 487506 285168 491234
rect 286428 487506 286456 491234
rect 287716 487506 287744 491234
rect 289004 487506 289032 491234
rect 290292 487506 290320 491234
rect 291580 487506 291608 491234
rect 274436 487478 274588 487506
rect 275724 487478 275968 487506
rect 277012 487478 277164 487506
rect 278392 487478 278728 487506
rect 279680 487478 280108 487506
rect 280968 487478 281396 487506
rect 282256 487478 282684 487506
rect 283544 487478 283972 487506
rect 284832 487478 285168 487506
rect 286120 487478 286456 487506
rect 287408 487478 287744 487506
rect 288696 487478 289032 487506
rect 289984 487478 290320 487506
rect 291272 487478 291608 487506
rect 292408 487506 292436 683198
rect 292500 491298 292528 696934
rect 292488 491292 292540 491298
rect 292488 491234 292540 491240
rect 293880 487778 293908 700703
rect 298008 700664 298060 700670
rect 298008 700606 298060 700612
rect 295248 700460 295300 700466
rect 295248 700402 295300 700408
rect 293834 487750 293908 487778
rect 292408 487478 292560 487506
rect 293834 487492 293862 487750
rect 295260 487506 295288 700402
rect 296628 700392 296680 700398
rect 296628 700334 296680 700340
rect 296640 487506 296668 700334
rect 298020 487506 298048 700606
rect 299400 487506 299428 700810
rect 300136 699718 300164 703520
rect 316040 701004 316092 701010
rect 316040 700946 316092 700952
rect 312544 700936 312596 700942
rect 312544 700878 312596 700884
rect 300768 700800 300820 700806
rect 300768 700742 300820 700748
rect 300124 699712 300176 699718
rect 300124 699654 300176 699660
rect 300780 487506 300808 700742
rect 302148 700256 302200 700262
rect 302148 700198 302200 700204
rect 302160 489914 302188 700198
rect 304908 700120 304960 700126
rect 304908 700062 304960 700068
rect 303528 700052 303580 700058
rect 303528 699994 303580 700000
rect 303540 489914 303568 699994
rect 304920 489914 304948 700062
rect 311992 699984 312044 699990
rect 311992 699926 312044 699932
rect 306288 699916 306340 699922
rect 306288 699858 306340 699864
rect 306300 491298 306328 699858
rect 310520 699848 310572 699854
rect 310520 699790 310572 699796
rect 307668 699780 307720 699786
rect 307668 699722 307720 699728
rect 307680 491298 307708 699722
rect 309140 699712 309192 699718
rect 309140 699654 309192 699660
rect 305828 491292 305880 491298
rect 305828 491234 305880 491240
rect 306288 491292 306340 491298
rect 306288 491234 306340 491240
rect 307116 491292 307168 491298
rect 307116 491234 307168 491240
rect 307668 491292 307720 491298
rect 307668 491234 307720 491240
rect 302068 489886 302188 489914
rect 303356 489886 303568 489914
rect 304644 489886 304948 489914
rect 302068 487506 302096 489886
rect 303356 487506 303384 489886
rect 304644 487506 304672 489886
rect 305840 487506 305868 491234
rect 307128 487506 307156 491234
rect 308404 491156 308456 491162
rect 308404 491098 308456 491104
rect 308416 487506 308444 491098
rect 295136 487478 295288 487506
rect 296424 487478 296668 487506
rect 297712 487478 298048 487506
rect 299092 487478 299428 487506
rect 300380 487478 300808 487506
rect 301668 487478 302096 487506
rect 302956 487478 303384 487506
rect 304244 487478 304672 487506
rect 305532 487478 305868 487506
rect 306820 487478 307156 487506
rect 308108 487478 308444 487506
rect 309152 487506 309180 699654
rect 310532 487506 310560 699790
rect 311900 491224 311952 491230
rect 311900 491166 311952 491172
rect 311912 487506 311940 491166
rect 312004 489914 312032 699926
rect 312556 491230 312584 700878
rect 315304 700528 315356 700534
rect 315304 700470 315356 700476
rect 313280 700188 313332 700194
rect 313280 700130 313332 700136
rect 313292 499574 313320 700130
rect 313292 499546 314148 499574
rect 312544 491224 312596 491230
rect 312544 491166 312596 491172
rect 312004 489886 312860 489914
rect 312832 487506 312860 489886
rect 314120 487506 314148 499546
rect 315316 491094 315344 700470
rect 316052 499574 316080 700946
rect 317420 700732 317472 700738
rect 317420 700674 317472 700680
rect 317432 499574 317460 700674
rect 324318 700632 324374 700641
rect 320180 700596 320232 700602
rect 324318 700567 324374 700576
rect 320180 700538 320232 700544
rect 319442 700496 319498 700505
rect 319442 700431 319498 700440
rect 316052 499546 316724 499574
rect 317432 499546 318012 499574
rect 315212 491088 315264 491094
rect 315212 491030 315264 491036
rect 315304 491088 315356 491094
rect 315304 491030 315356 491036
rect 315224 489914 315252 491030
rect 315224 489886 315436 489914
rect 315408 487506 315436 489886
rect 316696 487506 316724 499546
rect 317984 487506 318012 499546
rect 319456 491230 319484 700431
rect 320192 499574 320220 700538
rect 321560 700324 321612 700330
rect 321560 700266 321612 700272
rect 321572 499574 321600 700266
rect 323584 670744 323636 670750
rect 323584 670686 323636 670692
rect 320192 499546 320680 499574
rect 321572 499546 321968 499574
rect 319352 491224 319404 491230
rect 319352 491166 319404 491172
rect 319444 491224 319496 491230
rect 319444 491166 319496 491172
rect 319364 487506 319392 491166
rect 320652 487506 320680 499546
rect 321940 487506 321968 499546
rect 323596 491094 323624 670686
rect 324332 499574 324360 700567
rect 325698 700360 325754 700369
rect 325698 700295 325754 700304
rect 325712 499574 325740 700295
rect 332520 699786 332548 703520
rect 348804 702434 348832 703520
rect 347792 702406 348832 702434
rect 332508 699780 332560 699786
rect 332508 699722 332560 699728
rect 328460 683188 328512 683194
rect 328460 683130 328512 683136
rect 327724 618316 327776 618322
rect 327724 618258 327776 618264
rect 324332 499546 324544 499574
rect 325712 499546 325832 499574
rect 323308 491088 323360 491094
rect 323308 491030 323360 491036
rect 323584 491088 323636 491094
rect 323584 491030 323636 491036
rect 323320 487506 323348 491030
rect 324516 487506 324544 499546
rect 325804 487506 325832 499546
rect 327736 491298 327764 618258
rect 327724 491292 327776 491298
rect 327724 491234 327776 491240
rect 327172 491224 327224 491230
rect 327172 491166 327224 491172
rect 327184 487506 327212 491166
rect 328472 487506 328500 683130
rect 329840 656940 329892 656946
rect 329840 656882 329892 656888
rect 329852 487506 329880 656882
rect 332600 632120 332652 632126
rect 332600 632062 332652 632068
rect 331864 565888 331916 565894
rect 331864 565830 331916 565836
rect 331876 491230 331904 565830
rect 331864 491224 331916 491230
rect 331864 491166 331916 491172
rect 331220 491088 331272 491094
rect 331220 491030 331272 491036
rect 331232 487506 331260 491030
rect 332612 487506 332640 632062
rect 332692 605872 332744 605878
rect 332692 605814 332744 605820
rect 332704 499574 332732 605814
rect 335360 579692 335412 579698
rect 335360 579634 335412 579640
rect 334624 514820 334676 514826
rect 334624 514762 334676 514768
rect 332704 499546 333560 499574
rect 333532 487506 333560 499546
rect 334636 491094 334664 514762
rect 335372 499574 335400 579634
rect 336740 553444 336792 553450
rect 336740 553386 336792 553392
rect 336752 499574 336780 553386
rect 339500 527196 339552 527202
rect 339500 527138 339552 527144
rect 339512 499574 339540 527138
rect 340880 501016 340932 501022
rect 340880 500958 340932 500964
rect 340892 499574 340920 500958
rect 335372 499546 336136 499574
rect 336752 499546 337424 499574
rect 339512 499546 340000 499574
rect 340892 499546 341380 499574
rect 334900 491292 334952 491298
rect 334900 491234 334952 491240
rect 334624 491088 334676 491094
rect 334624 491030 334676 491036
rect 334912 487506 334940 491234
rect 336108 487506 336136 499546
rect 337396 487506 337424 499546
rect 338764 491224 338816 491230
rect 338764 491166 338816 491172
rect 338776 487506 338804 491166
rect 339972 487506 340000 499546
rect 341352 487506 341380 499546
rect 347792 491162 347820 702406
rect 364996 699922 365024 703520
rect 397472 700058 397500 703520
rect 413664 700126 413692 703520
rect 429856 700262 429884 703520
rect 462332 700874 462360 703520
rect 462320 700868 462372 700874
rect 462320 700810 462372 700816
rect 478524 700806 478552 703520
rect 478512 700800 478564 700806
rect 478512 700742 478564 700748
rect 494808 700670 494836 703520
rect 494796 700664 494848 700670
rect 494796 700606 494848 700612
rect 527192 700466 527220 703520
rect 527180 700460 527232 700466
rect 527180 700402 527232 700408
rect 543476 700398 543504 703520
rect 559668 700777 559696 703520
rect 559654 700768 559710 700777
rect 559654 700703 559710 700712
rect 543464 700392 543516 700398
rect 543464 700334 543516 700340
rect 429844 700256 429896 700262
rect 429844 700198 429896 700204
rect 413652 700120 413704 700126
rect 413652 700062 413704 700068
rect 397460 700052 397512 700058
rect 397460 699994 397512 700000
rect 364984 699916 365036 699922
rect 364984 699858 365036 699864
rect 580170 697232 580226 697241
rect 580170 697167 580226 697176
rect 580184 696998 580212 697167
rect 580172 696992 580224 696998
rect 580172 696934 580224 696940
rect 580170 683904 580226 683913
rect 580170 683839 580226 683848
rect 580184 683262 580212 683839
rect 580172 683256 580224 683262
rect 580172 683198 580224 683204
rect 580172 670812 580224 670818
rect 580172 670754 580224 670760
rect 580184 670721 580212 670754
rect 580170 670712 580226 670721
rect 580170 670647 580226 670656
rect 580170 644056 580226 644065
rect 580170 643991 580226 644000
rect 580184 643142 580212 643991
rect 580172 643136 580224 643142
rect 580172 643078 580224 643084
rect 580170 630864 580226 630873
rect 580170 630799 580226 630808
rect 580184 630698 580212 630799
rect 580172 630692 580224 630698
rect 580172 630634 580224 630640
rect 580170 617536 580226 617545
rect 580170 617471 580226 617480
rect 580184 616894 580212 617471
rect 580172 616888 580224 616894
rect 580172 616830 580224 616836
rect 579802 591016 579858 591025
rect 579802 590951 579858 590960
rect 579816 590714 579844 590951
rect 579804 590708 579856 590714
rect 579804 590650 579856 590656
rect 580170 577688 580226 577697
rect 580170 577623 580226 577632
rect 580184 576910 580212 577623
rect 580172 576904 580224 576910
rect 580172 576846 580224 576852
rect 579802 564360 579858 564369
rect 579802 564295 579858 564304
rect 579816 563106 579844 564295
rect 579804 563100 579856 563106
rect 579804 563042 579856 563048
rect 580170 537840 580226 537849
rect 580170 537775 580226 537784
rect 580184 536858 580212 537775
rect 580172 536852 580224 536858
rect 580172 536794 580224 536800
rect 580170 524512 580226 524521
rect 580170 524447 580172 524456
rect 580224 524447 580226 524456
rect 580172 524418 580224 524424
rect 580170 511320 580226 511329
rect 580170 511255 580226 511264
rect 580184 510678 580212 511255
rect 580172 510672 580224 510678
rect 580172 510614 580224 510620
rect 347780 491156 347832 491162
rect 347780 491098 347832 491104
rect 342720 491088 342772 491094
rect 342720 491030 342772 491036
rect 342732 487506 342760 491030
rect 385960 491020 386012 491026
rect 385960 490962 386012 490968
rect 346584 490884 346636 490890
rect 346584 490826 346636 490832
rect 344008 487620 344060 487626
rect 344008 487562 344060 487568
rect 345296 487620 345348 487626
rect 345296 487562 345348 487568
rect 344020 487506 344048 487562
rect 345308 487506 345336 487562
rect 346596 487506 346624 490826
rect 347964 490816 348016 490822
rect 347964 490758 348016 490764
rect 347976 487506 348004 490758
rect 349160 490748 349212 490754
rect 349160 490690 349212 490696
rect 349172 487506 349200 490690
rect 351920 490680 351972 490686
rect 351920 490622 351972 490628
rect 350540 490612 350592 490618
rect 350540 490554 350592 490560
rect 350552 487506 350580 490554
rect 351932 487506 351960 490622
rect 354312 490544 354364 490550
rect 354312 490486 354364 490492
rect 353300 490476 353352 490482
rect 353300 490418 353352 490424
rect 353312 487506 353340 490418
rect 354324 487506 354352 490486
rect 356888 490408 356940 490414
rect 356888 490350 356940 490356
rect 355600 487552 355652 487558
rect 309152 487478 309396 487506
rect 310532 487478 310684 487506
rect 311912 487478 311972 487506
rect 312832 487478 313260 487506
rect 314120 487478 314548 487506
rect 315408 487478 315836 487506
rect 316696 487478 317124 487506
rect 317984 487478 318412 487506
rect 319364 487478 319700 487506
rect 320652 487478 321080 487506
rect 321940 487478 322368 487506
rect 323320 487478 323656 487506
rect 324516 487478 324944 487506
rect 325804 487478 326232 487506
rect 327184 487478 327520 487506
rect 328472 487478 328808 487506
rect 329852 487478 330096 487506
rect 331232 487478 331384 487506
rect 332612 487478 332672 487506
rect 333532 487478 333960 487506
rect 334912 487478 335248 487506
rect 336108 487478 336536 487506
rect 337396 487478 337824 487506
rect 338776 487478 339112 487506
rect 339972 487478 340400 487506
rect 341352 487478 341780 487506
rect 342732 487478 343068 487506
rect 344020 487478 344356 487506
rect 345308 487478 345644 487506
rect 346596 487478 346932 487506
rect 347976 487478 348220 487506
rect 349172 487478 349508 487506
rect 350552 487478 350796 487506
rect 351932 487478 352084 487506
rect 353312 487478 353372 487506
rect 354324 487478 354660 487506
rect 356900 487506 356928 490350
rect 358176 490340 358228 490346
rect 358176 490282 358228 490288
rect 358188 487506 358216 490282
rect 360752 490272 360804 490278
rect 360752 490214 360804 490220
rect 385682 490240 385738 490249
rect 359464 487552 359516 487558
rect 355652 487500 355948 487506
rect 355600 487494 355948 487500
rect 355612 487478 355948 487494
rect 356900 487478 357236 487506
rect 358188 487478 358524 487506
rect 360764 487506 360792 490214
rect 362132 490204 362184 490210
rect 385682 490175 385738 490184
rect 362132 490146 362184 490152
rect 362144 487506 362172 490146
rect 364708 490136 364760 490142
rect 364708 490078 364760 490084
rect 384302 490104 384358 490113
rect 363420 487552 363472 487558
rect 359516 487500 359812 487506
rect 359464 487494 359812 487500
rect 359476 487478 359812 487494
rect 360764 487478 361100 487506
rect 362144 487478 362480 487506
rect 364720 487506 364748 490078
rect 365996 490068 366048 490074
rect 384302 490039 384358 490048
rect 365996 490010 366048 490016
rect 366008 487506 366036 490010
rect 368572 490000 368624 490006
rect 368572 489942 368624 489948
rect 367284 487552 367336 487558
rect 363472 487500 363768 487506
rect 363420 487494 363768 487500
rect 363432 487478 363768 487494
rect 364720 487478 365056 487506
rect 366008 487478 366344 487506
rect 368584 487506 368612 489942
rect 369860 489932 369912 489938
rect 369860 489874 369912 489880
rect 369872 487506 369900 489874
rect 384120 488504 384172 488510
rect 384120 488446 384172 488452
rect 383200 488436 383252 488442
rect 383200 488378 383252 488384
rect 383108 488164 383160 488170
rect 383108 488106 383160 488112
rect 383016 488028 383068 488034
rect 383016 487970 383068 487976
rect 382924 487892 382976 487898
rect 382924 487834 382976 487840
rect 371240 487620 371292 487626
rect 371240 487562 371292 487568
rect 371252 487506 371280 487562
rect 376300 487552 376352 487558
rect 367336 487500 367632 487506
rect 367284 487494 367632 487500
rect 367296 487478 367632 487494
rect 368584 487478 368920 487506
rect 369872 487478 370208 487506
rect 371252 487478 371496 487506
rect 376352 487500 376648 487506
rect 376300 487494 376648 487500
rect 376312 487478 376648 487494
rect 375012 487416 375064 487422
rect 375064 487364 375360 487370
rect 375012 487358 375360 487364
rect 375024 487342 375360 487358
rect 380176 487354 380512 487370
rect 380164 487348 380512 487354
rect 380216 487342 380512 487348
rect 380164 487290 380216 487296
rect 381452 487280 381504 487286
rect 378888 487218 379224 487234
rect 381504 487228 381800 487234
rect 381452 487222 381800 487228
rect 378876 487212 379224 487218
rect 378928 487206 379224 487212
rect 381464 487206 381800 487222
rect 378876 487154 378928 487160
rect 270868 487144 270920 487150
rect 240856 487082 241192 487098
rect 257692 487082 257936 487098
rect 258980 487082 259316 487098
rect 262844 487082 263180 487098
rect 266708 487082 267044 487098
rect 270572 487092 270868 487098
rect 270572 487086 270920 487092
rect 373906 487112 373962 487121
rect 240856 487076 241204 487082
rect 240856 487070 241152 487076
rect 257692 487076 257948 487082
rect 257692 487070 257896 487076
rect 241152 487018 241204 487024
rect 258980 487076 259328 487082
rect 258980 487070 259276 487076
rect 257896 487018 257948 487024
rect 262844 487076 263192 487082
rect 262844 487070 263140 487076
rect 259276 487018 259328 487024
rect 266708 487076 267056 487082
rect 266708 487070 267004 487076
rect 263140 487018 263192 487024
rect 270572 487070 270908 487086
rect 373906 487047 373962 487056
rect 267004 487018 267056 487024
rect 246304 487008 246356 487014
rect 246008 486956 246304 486962
rect 251272 487008 251324 487014
rect 246008 486950 246356 486956
rect 251160 486956 251272 486962
rect 252560 487008 252612 487014
rect 251160 486950 251324 486956
rect 252448 486956 252560 486962
rect 253848 487008 253900 487014
rect 252448 486950 252612 486956
rect 253736 486956 253848 486962
rect 256608 487008 256660 487014
rect 253736 486950 253900 486956
rect 256312 486956 256608 486962
rect 260564 487008 260616 487014
rect 256312 486950 256660 486956
rect 260268 486956 260564 486962
rect 261852 487008 261904 487014
rect 260268 486950 260616 486956
rect 261556 486956 261852 486962
rect 264428 487008 264480 487014
rect 261556 486950 261904 486956
rect 264132 486956 264428 486962
rect 265716 487008 265768 487014
rect 264132 486950 264480 486956
rect 265420 486956 265716 486962
rect 265420 486950 265768 486956
rect 372618 486976 372674 486985
rect 246008 486934 246344 486950
rect 251160 486934 251312 486950
rect 252448 486934 252600 486950
rect 253736 486934 253888 486950
rect 256312 486934 256648 486950
rect 260268 486934 260604 486950
rect 261556 486934 261892 486950
rect 264132 486934 264468 486950
rect 265420 486934 265756 486950
rect 373920 486962 373948 487047
rect 377586 486976 377642 486985
rect 372674 486934 372784 486962
rect 373920 486934 374072 486962
rect 372618 486911 372674 486920
rect 377642 486934 377936 486962
rect 377586 486911 377642 486920
rect 8022 486160 8078 486169
rect 8022 486095 8078 486104
rect 7932 462732 7984 462738
rect 7932 462674 7984 462680
rect 8036 97918 8064 486095
rect 234632 338014 235152 338042
rect 235276 338014 235428 338042
rect 235552 338014 235704 338042
rect 235828 338014 235980 338042
rect 236104 338014 236348 338042
rect 236472 338014 236624 338042
rect 236748 338014 236900 338042
rect 237024 338014 237176 338042
rect 237392 338014 237544 338042
rect 237668 338014 237820 338042
rect 237944 338014 238096 338042
rect 238220 338014 238372 338042
rect 238496 338014 238740 338042
rect 75828 336728 75880 336734
rect 75828 336670 75880 336676
rect 68928 336660 68980 336666
rect 68928 336602 68980 336608
rect 62028 336592 62080 336598
rect 62028 336534 62080 336540
rect 53748 336524 53800 336530
rect 53748 336466 53800 336472
rect 42708 336456 42760 336462
rect 42708 336398 42760 336404
rect 37188 336388 37240 336394
rect 37188 336330 37240 336336
rect 12346 336288 12402 336297
rect 12346 336223 12402 336232
rect 35808 336252 35860 336258
rect 10966 336152 11022 336161
rect 10966 336087 11022 336096
rect 8024 97912 8076 97918
rect 8024 97854 8076 97860
rect 7840 59356 7892 59362
rect 7840 59298 7892 59304
rect 7748 45552 7800 45558
rect 7748 45494 7800 45500
rect 7656 20188 7708 20194
rect 7656 20130 7708 20136
rect 8758 7576 8814 7585
rect 8758 7511 8814 7520
rect 7564 6656 7616 6662
rect 7564 6598 7616 6604
rect 7656 4956 7708 4962
rect 7656 4898 7708 4904
rect 6458 3360 6514 3369
rect 6458 3295 6514 3304
rect 6472 480 6500 3295
rect 7668 480 7696 4898
rect 8772 480 8800 7511
rect 10980 3534 11008 336087
rect 12254 7712 12310 7721
rect 12254 7647 12310 7656
rect 11152 3596 11204 3602
rect 11152 3538 11204 3544
rect 9956 3528 10008 3534
rect 9956 3470 10008 3476
rect 10968 3528 11020 3534
rect 10968 3470 11020 3476
rect 9968 480 9996 3470
rect 11164 480 11192 3538
rect 12268 3482 12296 7647
rect 12360 3602 12388 336223
rect 35808 336194 35860 336200
rect 28908 336184 28960 336190
rect 28908 336126 28960 336132
rect 19248 336116 19300 336122
rect 19248 336058 19300 336064
rect 13542 10296 13598 10305
rect 13542 10231 13598 10240
rect 12348 3596 12400 3602
rect 12348 3538 12400 3544
rect 12268 3454 12388 3482
rect 12360 480 12388 3454
rect 13556 480 13584 10231
rect 17038 7848 17094 7857
rect 17038 7783 17094 7792
rect 14738 3632 14794 3641
rect 14738 3567 14794 3576
rect 14752 480 14780 3567
rect 15934 3496 15990 3505
rect 15934 3431 15990 3440
rect 15948 480 15976 3431
rect 17052 480 17080 7783
rect 19260 3534 19288 336058
rect 20628 336048 20680 336054
rect 20628 335990 20680 335996
rect 19430 3768 19486 3777
rect 19430 3703 19486 3712
rect 18236 3528 18288 3534
rect 18236 3470 18288 3476
rect 19248 3528 19300 3534
rect 19248 3470 19300 3476
rect 18248 480 18276 3470
rect 19444 480 19472 3703
rect 20640 480 20668 335990
rect 26514 8936 26570 8945
rect 26514 8871 26570 8880
rect 21822 7984 21878 7993
rect 21822 7919 21878 7928
rect 21836 480 21864 7919
rect 25320 3596 25372 3602
rect 25320 3538 25372 3544
rect 24216 3528 24268 3534
rect 24216 3470 24268 3476
rect 23020 3460 23072 3466
rect 23020 3402 23072 3408
rect 23032 480 23060 3402
rect 24228 480 24256 3470
rect 25332 480 25360 3538
rect 26528 480 26556 8871
rect 28816 3664 28868 3670
rect 28816 3606 28868 3612
rect 27712 3392 27764 3398
rect 27712 3334 27764 3340
rect 27724 480 27752 3334
rect 28828 1850 28856 3606
rect 28920 3398 28948 336126
rect 30102 9072 30158 9081
rect 30102 9007 30158 9016
rect 28908 3392 28960 3398
rect 28908 3334 28960 3340
rect 28828 1822 28948 1850
rect 28920 480 28948 1822
rect 30116 480 30144 9007
rect 33600 8968 33652 8974
rect 33600 8910 33652 8916
rect 31300 3800 31352 3806
rect 31300 3742 31352 3748
rect 31312 480 31340 3742
rect 32404 3732 32456 3738
rect 32404 3674 32456 3680
rect 32416 480 32444 3674
rect 33612 480 33640 8910
rect 35820 3398 35848 336194
rect 37002 10432 37058 10441
rect 37002 10367 37058 10376
rect 35992 3868 36044 3874
rect 35992 3810 36044 3816
rect 34796 3392 34848 3398
rect 34796 3334 34848 3340
rect 35808 3392 35860 3398
rect 35808 3334 35860 3340
rect 34808 480 34836 3334
rect 36004 480 36032 3810
rect 37016 3482 37044 10367
rect 37200 6914 37228 336330
rect 41326 10568 41382 10577
rect 41326 10503 41382 10512
rect 37108 6886 37228 6914
rect 37108 3874 37136 6886
rect 39580 3936 39632 3942
rect 39580 3878 39632 3884
rect 37096 3868 37148 3874
rect 37096 3810 37148 3816
rect 38384 3868 38436 3874
rect 38384 3810 38436 3816
rect 37016 3454 37228 3482
rect 37200 480 37228 3454
rect 38396 480 38424 3810
rect 39592 480 39620 3878
rect 41340 3398 41368 10503
rect 42720 3398 42748 336398
rect 44088 336320 44140 336326
rect 44088 336262 44140 336268
rect 44100 3398 44128 336262
rect 45466 10704 45522 10713
rect 45466 10639 45522 10648
rect 45376 4004 45428 4010
rect 45376 3946 45428 3952
rect 40684 3392 40736 3398
rect 40684 3334 40736 3340
rect 41328 3392 41380 3398
rect 41328 3334 41380 3340
rect 41880 3392 41932 3398
rect 41880 3334 41932 3340
rect 42708 3392 42760 3398
rect 42708 3334 42760 3340
rect 43076 3392 43128 3398
rect 43076 3334 43128 3340
rect 44088 3392 44140 3398
rect 44088 3334 44140 3340
rect 44272 3392 44324 3398
rect 44272 3334 44324 3340
rect 40696 480 40724 3334
rect 41892 480 41920 3334
rect 43088 480 43116 3334
rect 44284 480 44312 3334
rect 45388 1986 45416 3946
rect 45480 3398 45508 10639
rect 53656 10396 53708 10402
rect 53656 10338 53708 10344
rect 49608 10328 49660 10334
rect 49608 10270 49660 10276
rect 47858 6216 47914 6225
rect 47858 6151 47914 6160
rect 46664 4072 46716 4078
rect 46664 4014 46716 4020
rect 45468 3392 45520 3398
rect 45468 3334 45520 3340
rect 45388 1958 45508 1986
rect 45480 480 45508 1958
rect 46676 480 46704 4014
rect 47872 480 47900 6151
rect 49620 3398 49648 10270
rect 51354 6352 51410 6361
rect 51354 6287 51410 6296
rect 50160 4140 50212 4146
rect 50160 4082 50212 4088
rect 48964 3392 49016 3398
rect 48964 3334 49016 3340
rect 49608 3392 49660 3398
rect 49608 3334 49660 3340
rect 48976 480 49004 3334
rect 50172 480 50200 4082
rect 51368 480 51396 6287
rect 53668 3398 53696 10338
rect 52552 3392 52604 3398
rect 52552 3334 52604 3340
rect 53656 3392 53708 3398
rect 53656 3334 53708 3340
rect 52564 480 52592 3334
rect 53760 480 53788 336466
rect 60648 10532 60700 10538
rect 60648 10474 60700 10480
rect 56508 10464 56560 10470
rect 56508 10406 56560 10412
rect 54942 6488 54998 6497
rect 54942 6423 54998 6432
rect 54956 480 54984 6423
rect 56520 3398 56548 10406
rect 58438 6624 58494 6633
rect 58438 6559 58494 6568
rect 56048 3392 56100 3398
rect 56048 3334 56100 3340
rect 56508 3392 56560 3398
rect 56508 3334 56560 3340
rect 56060 480 56088 3334
rect 57244 3324 57296 3330
rect 57244 3266 57296 3272
rect 57256 480 57284 3266
rect 58452 480 58480 6559
rect 60660 3398 60688 10474
rect 61936 6248 61988 6254
rect 61936 6190 61988 6196
rect 59636 3392 59688 3398
rect 59636 3334 59688 3340
rect 60648 3392 60700 3398
rect 60648 3334 60700 3340
rect 60832 3392 60884 3398
rect 60832 3334 60884 3340
rect 59648 480 59676 3334
rect 60844 480 60872 3334
rect 61948 3210 61976 6190
rect 62040 3398 62068 336534
rect 67548 10668 67600 10674
rect 67548 10610 67600 10616
rect 63224 10600 63276 10606
rect 63224 10542 63276 10548
rect 62028 3392 62080 3398
rect 62028 3334 62080 3340
rect 61948 3182 62068 3210
rect 62040 480 62068 3182
rect 63236 480 63264 10542
rect 65524 7608 65576 7614
rect 65524 7550 65576 7556
rect 64328 3256 64380 3262
rect 64328 3198 64380 3204
rect 64340 480 64368 3198
rect 65536 480 65564 7550
rect 67560 3398 67588 10610
rect 68940 3398 68968 336602
rect 74448 10804 74500 10810
rect 74448 10746 74500 10752
rect 70308 10736 70360 10742
rect 70308 10678 70360 10684
rect 69112 7676 69164 7682
rect 69112 7618 69164 7624
rect 66720 3392 66772 3398
rect 66720 3334 66772 3340
rect 67548 3392 67600 3398
rect 67548 3334 67600 3340
rect 67916 3392 67968 3398
rect 67916 3334 67968 3340
rect 68928 3392 68980 3398
rect 68928 3334 68980 3340
rect 66732 480 66760 3334
rect 67928 480 67956 3334
rect 69124 480 69152 7618
rect 70320 480 70348 10678
rect 72608 7744 72660 7750
rect 72608 7686 72660 7692
rect 71504 3188 71556 3194
rect 71504 3130 71556 3136
rect 71516 480 71544 3130
rect 72620 480 72648 7686
rect 74460 3262 74488 10746
rect 75840 3262 75868 336670
rect 82728 335980 82780 335986
rect 82728 335922 82780 335928
rect 79690 12064 79746 12073
rect 79690 11999 79746 12008
rect 78586 11792 78642 11801
rect 78586 11727 78642 11736
rect 76196 7812 76248 7818
rect 76196 7754 76248 7760
rect 73804 3256 73856 3262
rect 73804 3198 73856 3204
rect 74448 3256 74500 3262
rect 74448 3198 74500 3204
rect 75000 3256 75052 3262
rect 75000 3198 75052 3204
rect 75828 3256 75880 3262
rect 75828 3198 75880 3204
rect 73816 480 73844 3198
rect 75012 480 75040 3198
rect 76208 480 76236 7754
rect 78600 3262 78628 11727
rect 77392 3256 77444 3262
rect 77392 3198 77444 3204
rect 78588 3256 78640 3262
rect 78588 3198 78640 3204
rect 77404 480 77432 3198
rect 78588 3052 78640 3058
rect 78588 2994 78640 3000
rect 78600 480 78628 2994
rect 79704 480 79732 11999
rect 81346 11928 81402 11937
rect 81346 11863 81402 11872
rect 81360 3262 81388 11863
rect 82740 3262 82768 335922
rect 93768 335912 93820 335918
rect 93768 335854 93820 335860
rect 86868 335844 86920 335850
rect 86868 335786 86920 335792
rect 85488 11756 85540 11762
rect 85488 11698 85540 11704
rect 84108 10872 84160 10878
rect 84108 10814 84160 10820
rect 80888 3256 80940 3262
rect 80888 3198 80940 3204
rect 81348 3256 81400 3262
rect 81348 3198 81400 3204
rect 82084 3256 82136 3262
rect 82084 3198 82136 3204
rect 82728 3256 82780 3262
rect 82728 3198 82780 3204
rect 80900 480 80928 3198
rect 82096 480 82124 3198
rect 84120 3126 84148 10814
rect 85500 3262 85528 11698
rect 86684 10940 86736 10946
rect 86684 10882 86736 10888
rect 84476 3256 84528 3262
rect 84476 3198 84528 3204
rect 85488 3256 85540 3262
rect 85488 3198 85540 3204
rect 85672 3256 85724 3262
rect 85672 3198 85724 3204
rect 83280 3120 83332 3126
rect 83280 3062 83332 3068
rect 84108 3120 84160 3126
rect 84108 3062 84160 3068
rect 83292 480 83320 3062
rect 84488 480 84516 3198
rect 85684 480 85712 3198
rect 86696 3108 86724 10882
rect 86880 6914 86908 335786
rect 92388 11892 92440 11898
rect 92388 11834 92440 11840
rect 87972 11824 88024 11830
rect 87972 11766 88024 11772
rect 86788 6886 86908 6914
rect 86788 3262 86816 6886
rect 86776 3256 86828 3262
rect 86776 3198 86828 3204
rect 86696 3080 86908 3108
rect 86880 480 86908 3080
rect 87984 480 88012 11766
rect 91008 11008 91060 11014
rect 91008 10950 91060 10956
rect 91020 3262 91048 10950
rect 92400 3262 92428 11834
rect 90364 3256 90416 3262
rect 90364 3198 90416 3204
rect 91008 3256 91060 3262
rect 91008 3198 91060 3204
rect 91560 3256 91612 3262
rect 91560 3198 91612 3204
rect 92388 3256 92440 3262
rect 92388 3198 92440 3204
rect 89168 2984 89220 2990
rect 89168 2926 89220 2932
rect 89180 480 89208 2926
rect 90376 480 90404 3198
rect 91572 480 91600 3198
rect 93780 3126 93808 335854
rect 100668 335776 100720 335782
rect 100668 335718 100720 335724
rect 99288 13116 99340 13122
rect 99288 13058 99340 13064
rect 95148 11960 95200 11966
rect 95148 11902 95200 11908
rect 95056 10260 95108 10266
rect 95056 10202 95108 10208
rect 95068 3126 95096 10202
rect 92756 3120 92808 3126
rect 92756 3062 92808 3068
rect 93768 3120 93820 3126
rect 93768 3062 93820 3068
rect 93952 3120 94004 3126
rect 93952 3062 94004 3068
rect 95056 3120 95108 3126
rect 95056 3062 95108 3068
rect 92768 480 92796 3062
rect 93964 480 93992 3062
rect 95160 480 95188 11902
rect 97908 10192 97960 10198
rect 97908 10134 97960 10140
rect 97920 3126 97948 10134
rect 99300 3126 99328 13058
rect 100680 3126 100708 335718
rect 107568 335708 107620 335714
rect 107568 335650 107620 335656
rect 106188 13252 106240 13258
rect 106188 13194 106240 13200
rect 103428 13184 103480 13190
rect 103428 13126 103480 13132
rect 102048 10124 102100 10130
rect 102048 10066 102100 10072
rect 97448 3120 97500 3126
rect 97448 3062 97500 3068
rect 97908 3120 97960 3126
rect 97908 3062 97960 3068
rect 98644 3120 98696 3126
rect 98644 3062 98696 3068
rect 99288 3120 99340 3126
rect 99288 3062 99340 3068
rect 99840 3120 99892 3126
rect 99840 3062 99892 3068
rect 100668 3120 100720 3126
rect 100668 3062 100720 3068
rect 96252 2984 96304 2990
rect 96252 2926 96304 2932
rect 96264 480 96292 2926
rect 97460 480 97488 3062
rect 98656 480 98684 3062
rect 99852 480 99880 3062
rect 102060 2922 102088 10066
rect 103440 2990 103468 13126
rect 104532 10056 104584 10062
rect 104532 9998 104584 10004
rect 102232 2984 102284 2990
rect 102232 2926 102284 2932
rect 103428 2984 103480 2990
rect 103428 2926 103480 2932
rect 101036 2916 101088 2922
rect 101036 2858 101088 2864
rect 102048 2916 102100 2922
rect 102048 2858 102100 2864
rect 101048 480 101076 2858
rect 102244 480 102272 2926
rect 103336 2916 103388 2922
rect 103336 2858 103388 2864
rect 103348 480 103376 2858
rect 104544 480 104572 9998
rect 106200 2990 106228 13194
rect 107580 2990 107608 335650
rect 114468 335640 114520 335646
rect 114468 335582 114520 335588
rect 112812 13388 112864 13394
rect 112812 13330 112864 13336
rect 110328 13320 110380 13326
rect 110328 13262 110380 13268
rect 108948 9988 109000 9994
rect 108948 9930 109000 9936
rect 108960 2990 108988 9930
rect 110340 2990 110368 13262
rect 111616 9920 111668 9926
rect 111616 9862 111668 9868
rect 105728 2984 105780 2990
rect 105728 2926 105780 2932
rect 106188 2984 106240 2990
rect 106188 2926 106240 2932
rect 106924 2984 106976 2990
rect 106924 2926 106976 2932
rect 107568 2984 107620 2990
rect 107568 2926 107620 2932
rect 108120 2984 108172 2990
rect 108120 2926 108172 2932
rect 108948 2984 109000 2990
rect 108948 2926 109000 2932
rect 109316 2984 109368 2990
rect 109316 2926 109368 2932
rect 110328 2984 110380 2990
rect 110328 2926 110380 2932
rect 105740 480 105768 2926
rect 106936 480 106964 2926
rect 108132 480 108160 2926
rect 109328 480 109356 2926
rect 110512 2916 110564 2922
rect 110512 2858 110564 2864
rect 110524 480 110552 2858
rect 111628 480 111656 9862
rect 112824 480 112852 13330
rect 114480 2854 114508 335582
rect 121368 335572 121420 335578
rect 121368 335514 121420 335520
rect 119896 13524 119948 13530
rect 119896 13466 119948 13472
rect 117228 13456 117280 13462
rect 117228 13398 117280 13404
rect 115848 9852 115900 9858
rect 115848 9794 115900 9800
rect 115860 2854 115888 9794
rect 117240 2854 117268 13398
rect 119804 9784 119856 9790
rect 119804 9726 119856 9732
rect 119816 2854 119844 9726
rect 114008 2848 114060 2854
rect 114008 2790 114060 2796
rect 114468 2848 114520 2854
rect 114468 2790 114520 2796
rect 115204 2848 115256 2854
rect 115204 2790 115256 2796
rect 115848 2848 115900 2854
rect 115848 2790 115900 2796
rect 116400 2848 116452 2854
rect 116400 2790 116452 2796
rect 117228 2848 117280 2854
rect 117228 2790 117280 2796
rect 117596 2848 117648 2854
rect 117596 2790 117648 2796
rect 118792 2848 118844 2854
rect 118792 2790 118844 2796
rect 119804 2848 119856 2854
rect 119804 2790 119856 2796
rect 114020 480 114048 2790
rect 115216 480 115244 2790
rect 116412 480 116440 2790
rect 117608 480 117636 2790
rect 118804 480 118832 2790
rect 119908 480 119936 13466
rect 121380 6914 121408 335514
rect 193864 335504 193916 335510
rect 193864 335446 193916 335452
rect 191104 335436 191156 335442
rect 191104 335378 191156 335384
rect 161296 12436 161348 12442
rect 161296 12378 161348 12384
rect 160100 12368 160152 12374
rect 160100 12310 160152 12316
rect 147588 12300 147640 12306
rect 147588 12242 147640 12248
rect 144828 12232 144880 12238
rect 144828 12174 144880 12180
rect 140044 12164 140096 12170
rect 140044 12106 140096 12112
rect 136456 12096 136508 12102
rect 136456 12038 136508 12044
rect 125876 12028 125928 12034
rect 125876 11970 125928 11976
rect 122748 9716 122800 9722
rect 122748 9658 122800 9664
rect 121104 6886 121408 6914
rect 121104 480 121132 6886
rect 122300 598 122512 626
rect 122300 480 122328 598
rect 122484 490 122512 598
rect 122760 490 122788 9658
rect 123484 5364 123536 5370
rect 123484 5306 123536 5312
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9926 -960 10038 480
rect 11122 -960 11234 480
rect 12318 -960 12430 480
rect 13514 -960 13626 480
rect 14710 -960 14822 480
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 18206 -960 18318 480
rect 19402 -960 19514 480
rect 20598 -960 20710 480
rect 21794 -960 21906 480
rect 22990 -960 23102 480
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26486 -960 26598 480
rect 27682 -960 27794 480
rect 28878 -960 28990 480
rect 30074 -960 30186 480
rect 31270 -960 31382 480
rect 32374 -960 32486 480
rect 33570 -960 33682 480
rect 34766 -960 34878 480
rect 35962 -960 36074 480
rect 37158 -960 37270 480
rect 38354 -960 38466 480
rect 39550 -960 39662 480
rect 40654 -960 40766 480
rect 41850 -960 41962 480
rect 43046 -960 43158 480
rect 44242 -960 44354 480
rect 45438 -960 45550 480
rect 46634 -960 46746 480
rect 47830 -960 47942 480
rect 48934 -960 49046 480
rect 50130 -960 50242 480
rect 51326 -960 51438 480
rect 52522 -960 52634 480
rect 53718 -960 53830 480
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 57214 -960 57326 480
rect 58410 -960 58522 480
rect 59606 -960 59718 480
rect 60802 -960 60914 480
rect 61998 -960 62110 480
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65494 -960 65606 480
rect 66690 -960 66802 480
rect 67886 -960 67998 480
rect 69082 -960 69194 480
rect 70278 -960 70390 480
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73774 -960 73886 480
rect 74970 -960 75082 480
rect 76166 -960 76278 480
rect 77362 -960 77474 480
rect 78558 -960 78670 480
rect 79662 -960 79774 480
rect 80858 -960 80970 480
rect 82054 -960 82166 480
rect 83250 -960 83362 480
rect 84446 -960 84558 480
rect 85642 -960 85754 480
rect 86838 -960 86950 480
rect 87942 -960 88054 480
rect 89138 -960 89250 480
rect 90334 -960 90446 480
rect 91530 -960 91642 480
rect 92726 -960 92838 480
rect 93922 -960 94034 480
rect 95118 -960 95230 480
rect 96222 -960 96334 480
rect 97418 -960 97530 480
rect 98614 -960 98726 480
rect 99810 -960 99922 480
rect 101006 -960 101118 480
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104502 -960 104614 480
rect 105698 -960 105810 480
rect 106894 -960 107006 480
rect 108090 -960 108202 480
rect 109286 -960 109398 480
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112782 -960 112894 480
rect 113978 -960 114090 480
rect 115174 -960 115286 480
rect 116370 -960 116482 480
rect 117566 -960 117678 480
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 121062 -960 121174 480
rect 122258 -960 122370 480
rect 122484 462 122788 490
rect 123496 480 123524 5306
rect 124680 5296 124732 5302
rect 124680 5238 124732 5244
rect 124692 480 124720 5238
rect 125888 480 125916 11970
rect 135258 9344 135314 9353
rect 135258 9279 135314 9288
rect 131762 9208 131818 9217
rect 131762 9143 131818 9152
rect 128176 7880 128228 7886
rect 128176 7822 128228 7828
rect 126980 6316 127032 6322
rect 126980 6258 127032 6264
rect 126992 480 127020 6258
rect 128188 480 128216 7822
rect 130568 6384 130620 6390
rect 130568 6326 130620 6332
rect 129370 4856 129426 4865
rect 129370 4791 129426 4800
rect 129384 480 129412 4791
rect 130580 480 130608 6326
rect 131776 480 131804 9143
rect 134156 7948 134208 7954
rect 134156 7890 134208 7896
rect 132958 4992 133014 5001
rect 132958 4927 133014 4936
rect 132972 480 133000 4927
rect 134168 480 134196 7890
rect 135272 480 135300 9279
rect 136468 480 136496 12038
rect 138848 9036 138900 9042
rect 138848 8978 138900 8984
rect 137652 8016 137704 8022
rect 137652 7958 137704 7964
rect 137664 480 137692 7958
rect 138860 480 138888 8978
rect 140056 480 140084 12106
rect 142436 9104 142488 9110
rect 142436 9046 142488 9052
rect 141240 8084 141292 8090
rect 141240 8026 141292 8032
rect 141252 480 141280 8026
rect 142448 480 142476 9046
rect 144736 8152 144788 8158
rect 144736 8094 144788 8100
rect 143540 4208 143592 4214
rect 143540 4150 143592 4156
rect 143552 480 143580 4150
rect 144748 480 144776 8094
rect 144840 4214 144868 12174
rect 145932 9172 145984 9178
rect 145932 9114 145984 9120
rect 144828 4208 144880 4214
rect 144828 4150 144880 4156
rect 145944 480 145972 9114
rect 147140 598 147352 626
rect 147140 480 147168 598
rect 147324 490 147352 598
rect 147600 490 147628 12242
rect 156604 9376 156656 9382
rect 156604 9318 156656 9324
rect 153016 9308 153068 9314
rect 153016 9250 153068 9256
rect 149520 9240 149572 9246
rect 149520 9182 149572 9188
rect 148324 8220 148376 8226
rect 148324 8162 148376 8168
rect 123454 -960 123566 480
rect 124650 -960 124762 480
rect 125846 -960 125958 480
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 129342 -960 129454 480
rect 130538 -960 130650 480
rect 131734 -960 131846 480
rect 132930 -960 133042 480
rect 134126 -960 134238 480
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137622 -960 137734 480
rect 138818 -960 138930 480
rect 140014 -960 140126 480
rect 141210 -960 141322 480
rect 142406 -960 142518 480
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145902 -960 146014 480
rect 147098 -960 147210 480
rect 147324 462 147628 490
rect 148336 480 148364 8162
rect 149532 480 149560 9182
rect 151820 8288 151872 8294
rect 151820 8230 151872 8236
rect 150624 6452 150676 6458
rect 150624 6394 150676 6400
rect 150636 480 150664 6394
rect 151832 480 151860 8230
rect 153028 480 153056 9250
rect 155408 7540 155460 7546
rect 155408 7482 155460 7488
rect 154212 6520 154264 6526
rect 154212 6462 154264 6468
rect 154224 480 154252 6462
rect 155420 480 155448 7482
rect 156616 480 156644 9318
rect 158904 7472 158956 7478
rect 158904 7414 158956 7420
rect 157800 6588 157852 6594
rect 157800 6530 157852 6536
rect 157812 480 157840 6530
rect 158916 480 158944 7414
rect 160112 480 160140 12310
rect 161308 480 161336 12378
rect 164884 11688 164936 11694
rect 164884 11630 164936 11636
rect 163688 7404 163740 7410
rect 163688 7346 163740 7352
rect 162492 6656 162544 6662
rect 162492 6598 162544 6604
rect 162504 480 162532 6598
rect 163700 480 163728 7346
rect 164896 480 164924 11630
rect 174268 11620 174320 11626
rect 174268 11562 174320 11568
rect 167184 7336 167236 7342
rect 167184 7278 167236 7284
rect 166080 6724 166132 6730
rect 166080 6666 166132 6672
rect 166092 480 166120 6666
rect 167196 480 167224 7278
rect 170772 7268 170824 7274
rect 170772 7210 170824 7216
rect 169576 6792 169628 6798
rect 169576 6734 169628 6740
rect 168378 5264 168434 5273
rect 168378 5199 168434 5208
rect 168392 480 168420 5199
rect 169588 480 169616 6734
rect 170784 480 170812 7210
rect 173164 6860 173216 6866
rect 173164 6802 173216 6808
rect 171968 4548 172020 4554
rect 171968 4490 172020 4496
rect 171980 480 172008 4490
rect 173176 480 173204 6802
rect 174280 480 174308 11562
rect 177856 11552 177908 11558
rect 177856 11494 177908 11500
rect 176660 6112 176712 6118
rect 176660 6054 176712 6060
rect 175462 5128 175518 5137
rect 175462 5063 175518 5072
rect 175476 480 175504 5063
rect 176672 480 176700 6054
rect 177868 480 177896 11494
rect 181444 11484 181496 11490
rect 181444 11426 181496 11432
rect 180248 6044 180300 6050
rect 180248 5986 180300 5992
rect 179052 5024 179104 5030
rect 179052 4966 179104 4972
rect 179064 480 179092 4966
rect 180260 480 180288 5986
rect 181456 480 181484 11426
rect 184940 11416 184992 11422
rect 184940 11358 184992 11364
rect 183744 5976 183796 5982
rect 183744 5918 183796 5924
rect 182548 5092 182600 5098
rect 182548 5034 182600 5040
rect 182560 480 182588 5034
rect 183756 480 183784 5918
rect 184952 480 184980 11358
rect 188528 9444 188580 9450
rect 188528 9386 188580 9392
rect 187332 5908 187384 5914
rect 187332 5850 187384 5856
rect 186136 5160 186188 5166
rect 186136 5102 186188 5108
rect 186148 480 186176 5102
rect 187344 480 187372 5850
rect 188540 480 188568 9386
rect 190828 5840 190880 5846
rect 190828 5782 190880 5788
rect 189724 5228 189776 5234
rect 189724 5170 189776 5176
rect 189736 480 189764 5170
rect 190840 480 190868 5782
rect 191116 5370 191144 335378
rect 192024 9512 192076 9518
rect 192024 9454 192076 9460
rect 191104 5364 191156 5370
rect 191104 5306 191156 5312
rect 192036 480 192064 9454
rect 193220 5364 193272 5370
rect 193220 5306 193272 5312
rect 193232 480 193260 5306
rect 193876 5302 193904 335446
rect 234632 11665 234660 338014
rect 235276 335354 235304 338014
rect 234816 335326 235304 335354
rect 234712 326392 234764 326398
rect 234712 326334 234764 326340
rect 234618 11656 234674 11665
rect 234618 11591 234674 11600
rect 205548 11348 205600 11354
rect 205548 11290 205600 11296
rect 199108 9648 199160 9654
rect 199108 9590 199160 9596
rect 195612 9580 195664 9586
rect 195612 9522 195664 9528
rect 194416 5772 194468 5778
rect 194416 5714 194468 5720
rect 193864 5296 193916 5302
rect 193864 5238 193916 5244
rect 194428 480 194456 5714
rect 195624 480 195652 9522
rect 197912 5704 197964 5710
rect 197912 5646 197964 5652
rect 196808 5364 196860 5370
rect 196808 5306 196860 5312
rect 196820 480 196848 5306
rect 197924 480 197952 5646
rect 199120 480 199148 9590
rect 202696 8900 202748 8906
rect 202696 8842 202748 8848
rect 201500 5636 201552 5642
rect 201500 5578 201552 5584
rect 200304 5432 200356 5438
rect 200304 5374 200356 5380
rect 200316 480 200344 5374
rect 201512 480 201540 5578
rect 202708 480 202736 8842
rect 203892 5500 203944 5506
rect 203892 5442 203944 5448
rect 203904 480 203932 5442
rect 205100 598 205312 626
rect 205100 480 205128 598
rect 205284 490 205312 598
rect 205560 490 205588 11290
rect 209044 11280 209096 11286
rect 209044 11222 209096 11228
rect 206192 8832 206244 8838
rect 206192 8774 206244 8780
rect 148294 -960 148406 480
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 154182 -960 154294 480
rect 155378 -960 155490 480
rect 156574 -960 156686 480
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162462 -960 162574 480
rect 163658 -960 163770 480
rect 164854 -960 164966 480
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170742 -960 170854 480
rect 171938 -960 172050 480
rect 173134 -960 173246 480
rect 174238 -960 174350 480
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 179022 -960 179134 480
rect 180218 -960 180330 480
rect 181414 -960 181526 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 187302 -960 187414 480
rect 188498 -960 188610 480
rect 189694 -960 189806 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 199078 -960 199190 480
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 205284 462 205588 490
rect 206204 480 206232 8774
rect 207388 4752 207440 4758
rect 207388 4694 207440 4700
rect 207400 480 207428 4694
rect 208596 598 208808 626
rect 208596 480 208624 598
rect 208780 490 208808 598
rect 209056 490 209084 11222
rect 212172 11212 212224 11218
rect 212172 11154 212224 11160
rect 209780 8764 209832 8770
rect 209780 8706 209832 8712
rect 206162 -960 206274 480
rect 207358 -960 207470 480
rect 208554 -960 208666 480
rect 208780 462 209084 490
rect 209792 480 209820 8706
rect 210976 4684 211028 4690
rect 210976 4626 211028 4632
rect 210988 480 211016 4626
rect 212184 480 212212 11154
rect 215668 11144 215720 11150
rect 215668 11086 215720 11092
rect 213368 8696 213420 8702
rect 213368 8638 213420 8644
rect 213380 480 213408 8638
rect 214472 4616 214524 4622
rect 214472 4558 214524 4564
rect 214484 480 214512 4558
rect 215680 480 215708 11086
rect 216864 8628 216916 8634
rect 216864 8570 216916 8576
rect 216876 480 216904 8570
rect 220452 8560 220504 8566
rect 220452 8502 220504 8508
rect 219256 6996 219308 7002
rect 219256 6938 219308 6944
rect 218060 4208 218112 4214
rect 218060 4150 218112 4156
rect 218072 480 218100 4150
rect 219268 480 219296 6938
rect 220464 480 220492 8502
rect 223948 8492 224000 8498
rect 223948 8434 224000 8440
rect 222752 7200 222804 7206
rect 222752 7142 222804 7148
rect 221556 4480 221608 4486
rect 221556 4422 221608 4428
rect 221568 480 221596 4422
rect 222764 480 222792 7142
rect 223960 480 223988 8434
rect 227536 8424 227588 8430
rect 227536 8366 227588 8372
rect 226340 5568 226392 5574
rect 226340 5510 226392 5516
rect 225144 4412 225196 4418
rect 225144 4354 225196 4360
rect 225156 480 225184 4354
rect 226352 480 226380 5510
rect 227548 480 227576 8366
rect 231032 8356 231084 8362
rect 231032 8298 231084 8304
rect 229836 7132 229888 7138
rect 229836 7074 229888 7080
rect 228732 4344 228784 4350
rect 228732 4286 228784 4292
rect 228744 480 228772 4286
rect 229848 480 229876 7074
rect 231044 480 231072 8298
rect 233424 7064 233476 7070
rect 233424 7006 233476 7012
rect 232228 4820 232280 4826
rect 232228 4762 232280 4768
rect 232240 480 232268 4762
rect 233436 480 233464 7006
rect 234620 4956 234672 4962
rect 234620 4898 234672 4904
rect 234632 480 234660 4898
rect 234724 4894 234752 326334
rect 234712 4888 234764 4894
rect 234712 4830 234764 4836
rect 234816 4282 234844 335326
rect 235552 326398 235580 338014
rect 235540 326392 235592 326398
rect 235540 326334 235592 326340
rect 235828 316034 235856 338014
rect 236104 336025 236132 338014
rect 236090 336016 236146 336025
rect 236090 335951 236146 335960
rect 236092 326392 236144 326398
rect 236092 326334 236144 326340
rect 234908 316006 235856 316034
rect 234908 6186 234936 316006
rect 234896 6180 234948 6186
rect 234896 6122 234948 6128
rect 236104 4894 236132 326334
rect 236184 323196 236236 323202
rect 236184 323138 236236 323144
rect 236196 7585 236224 323138
rect 236472 316034 236500 338014
rect 236748 326398 236776 338014
rect 236736 326392 236788 326398
rect 236736 326334 236788 326340
rect 237024 323202 237052 338014
rect 237392 336161 237420 338014
rect 237668 336297 237696 338014
rect 237654 336288 237710 336297
rect 237654 336223 237710 336232
rect 237378 336152 237434 336161
rect 237378 336087 237434 336096
rect 237944 335354 237972 338014
rect 237484 335326 237972 335354
rect 237380 326392 237432 326398
rect 237380 326334 237432 326340
rect 237012 323196 237064 323202
rect 237012 323138 237064 323144
rect 236288 316006 236500 316034
rect 236182 7576 236238 7585
rect 236182 7511 236238 7520
rect 236092 4888 236144 4894
rect 236092 4830 236144 4836
rect 234804 4276 234856 4282
rect 234804 4218 234856 4224
rect 235816 4276 235868 4282
rect 235816 4218 235868 4224
rect 235828 480 235856 4218
rect 236288 3369 236316 316006
rect 237012 4888 237064 4894
rect 237012 4830 237064 4836
rect 236274 3360 236330 3369
rect 236274 3295 236330 3304
rect 237024 480 237052 4830
rect 237392 3641 237420 326334
rect 237484 7721 237512 335326
rect 238220 316034 238248 338014
rect 238496 326398 238524 338014
rect 239002 337770 239030 338028
rect 239140 338014 239292 338042
rect 239416 338014 239568 338042
rect 239692 338014 239936 338042
rect 240152 338014 240212 338042
rect 240428 338014 240488 338042
rect 240612 338014 240764 338042
rect 240888 338014 241132 338042
rect 241256 338014 241408 338042
rect 239002 337742 239076 337770
rect 239048 328454 239076 337742
rect 238956 328426 239076 328454
rect 238484 326392 238536 326398
rect 238484 326334 238536 326340
rect 238852 326392 238904 326398
rect 238852 326334 238904 326340
rect 237576 316006 238248 316034
rect 237576 10305 237604 316006
rect 237562 10296 237618 10305
rect 237562 10231 237618 10240
rect 237470 7712 237526 7721
rect 237470 7647 237526 7656
rect 238116 6180 238168 6186
rect 238116 6122 238168 6128
rect 237378 3632 237434 3641
rect 237378 3567 237434 3576
rect 238128 480 238156 6122
rect 238864 3777 238892 326334
rect 238956 323626 238984 328426
rect 238956 323598 239076 323626
rect 238944 319592 238996 319598
rect 238944 319534 238996 319540
rect 238956 7857 238984 319534
rect 238942 7848 238998 7857
rect 238942 7783 238998 7792
rect 238850 3768 238906 3777
rect 238850 3703 238906 3712
rect 239048 3505 239076 323598
rect 239140 319598 239168 338014
rect 239416 336122 239444 338014
rect 239404 336116 239456 336122
rect 239404 336058 239456 336064
rect 239692 326398 239720 338014
rect 240152 336054 240180 338014
rect 240140 336048 240192 336054
rect 240140 335990 240192 335996
rect 239680 326392 239732 326398
rect 239680 326334 239732 326340
rect 240324 326392 240376 326398
rect 240324 326334 240376 326340
rect 240232 321904 240284 321910
rect 240232 321846 240284 321852
rect 239128 319592 239180 319598
rect 239128 319534 239180 319540
rect 239034 3496 239090 3505
rect 240244 3466 240272 321846
rect 240336 3534 240364 326334
rect 240428 7993 240456 338014
rect 240612 321910 240640 338014
rect 240888 326398 240916 338014
rect 240876 326392 240928 326398
rect 240876 326334 240928 326340
rect 240600 321904 240652 321910
rect 240600 321846 240652 321852
rect 241256 316034 241284 338014
rect 241670 337770 241698 338028
rect 241808 338014 241960 338042
rect 242084 338014 242328 338042
rect 242452 338014 242604 338042
rect 242728 338014 242880 338042
rect 243096 338014 243156 338042
rect 243280 338014 243524 338042
rect 243648 338014 243800 338042
rect 243924 338014 244076 338042
rect 244352 338014 244504 338042
rect 241670 337742 241744 337770
rect 241612 326392 241664 326398
rect 241612 326334 241664 326340
rect 240520 316006 241284 316034
rect 240414 7984 240470 7993
rect 240414 7919 240470 7928
rect 240520 3602 240548 316006
rect 241624 3670 241652 326334
rect 241716 8945 241744 337742
rect 241808 336190 241836 338014
rect 241796 336184 241848 336190
rect 241796 336126 241848 336132
rect 242084 326398 242112 338014
rect 242452 335354 242480 338014
rect 242176 335326 242480 335354
rect 242072 326392 242124 326398
rect 242072 326334 242124 326340
rect 242176 321554 242204 335326
rect 241808 321526 242204 321554
rect 241808 9081 241836 321526
rect 242728 316034 242756 338014
rect 243096 328454 243124 338014
rect 243280 335354 243308 338014
rect 243648 336258 243676 338014
rect 243924 336394 243952 338014
rect 243912 336388 243964 336394
rect 243912 336330 243964 336336
rect 243636 336252 243688 336258
rect 243636 336194 243688 336200
rect 243004 328426 243124 328454
rect 243188 335326 243308 335354
rect 243544 335368 243596 335374
rect 243004 323762 243032 328426
rect 243004 323734 243124 323762
rect 242992 323604 243044 323610
rect 242992 323546 243044 323552
rect 241900 316006 242756 316034
rect 241794 9072 241850 9081
rect 241794 9007 241850 9016
rect 241702 8936 241758 8945
rect 241702 8871 241758 8880
rect 241900 3806 241928 316006
rect 243004 8974 243032 323546
rect 242992 8968 243044 8974
rect 242992 8910 243044 8916
rect 241888 3800 241940 3806
rect 241888 3742 241940 3748
rect 243096 3738 243124 323734
rect 243188 323610 243216 335326
rect 243544 335310 243596 335316
rect 243176 323604 243228 323610
rect 243176 323546 243228 323552
rect 243556 5273 243584 335310
rect 244372 326392 244424 326398
rect 244372 326334 244424 326340
rect 243542 5264 243598 5273
rect 243542 5199 243598 5208
rect 244096 4072 244148 4078
rect 244096 4014 244148 4020
rect 243084 3732 243136 3738
rect 243084 3674 243136 3680
rect 241612 3664 241664 3670
rect 241612 3606 241664 3612
rect 241704 3664 241756 3670
rect 241704 3606 241756 3612
rect 240508 3596 240560 3602
rect 240508 3538 240560 3544
rect 240324 3528 240376 3534
rect 240324 3470 240376 3476
rect 240506 3496 240562 3505
rect 239034 3431 239090 3440
rect 240232 3460 240284 3466
rect 240506 3431 240562 3440
rect 240232 3402 240284 3408
rect 239310 3360 239366 3369
rect 239310 3295 239366 3304
rect 239324 480 239352 3295
rect 240520 480 240548 3431
rect 241716 480 241744 3606
rect 242900 3460 242952 3466
rect 242900 3402 242952 3408
rect 242912 480 242940 3402
rect 244108 480 244136 4014
rect 244384 3942 244412 326334
rect 244476 10441 244504 338014
rect 244660 338014 244720 338042
rect 244844 338014 244996 338042
rect 245120 338014 245272 338042
rect 245396 338014 245548 338042
rect 245672 338014 245916 338042
rect 246040 338014 246192 338042
rect 246316 338014 246468 338042
rect 246592 338014 246744 338042
rect 244556 326460 244608 326466
rect 244556 326402 244608 326408
rect 244568 10577 244596 326402
rect 244554 10568 244610 10577
rect 244554 10503 244610 10512
rect 244462 10432 244518 10441
rect 244462 10367 244518 10376
rect 244372 3936 244424 3942
rect 244372 3878 244424 3884
rect 244660 3874 244688 338014
rect 244844 326398 244872 338014
rect 245016 336388 245068 336394
rect 245016 336330 245068 336336
rect 244924 336184 244976 336190
rect 244924 336126 244976 336132
rect 244832 326392 244884 326398
rect 244832 326334 244884 326340
rect 244936 4826 244964 336126
rect 244924 4820 244976 4826
rect 244924 4762 244976 4768
rect 245028 4554 245056 336330
rect 245120 326466 245148 338014
rect 245396 336462 245424 338014
rect 245384 336456 245436 336462
rect 245384 336398 245436 336404
rect 245672 336326 245700 338014
rect 245660 336320 245712 336326
rect 245660 336262 245712 336268
rect 246040 335354 246068 338014
rect 245856 335326 246068 335354
rect 245108 326460 245160 326466
rect 245108 326402 245160 326408
rect 245752 326392 245804 326398
rect 245752 326334 245804 326340
rect 245016 4548 245068 4554
rect 245016 4490 245068 4496
rect 245764 4010 245792 326334
rect 245856 10713 245884 335326
rect 245936 326460 245988 326466
rect 245936 326402 245988 326408
rect 245842 10704 245898 10713
rect 245842 10639 245898 10648
rect 245948 4146 245976 326402
rect 246316 326398 246344 338014
rect 246396 336320 246448 336326
rect 246396 336262 246448 336268
rect 246304 326392 246356 326398
rect 246304 326334 246356 326340
rect 246408 316034 246436 336262
rect 246592 326466 246620 338014
rect 247098 337770 247126 338028
rect 247374 337770 247402 338028
rect 247512 338014 247664 338042
rect 247788 338014 247940 338042
rect 248064 338014 248308 338042
rect 248432 338014 248584 338042
rect 248708 338014 248860 338042
rect 248984 338014 249136 338042
rect 249260 338014 249504 338042
rect 249628 338014 249780 338042
rect 249996 338014 250056 338042
rect 250180 338014 250332 338042
rect 250456 338014 250700 338042
rect 250824 338014 250976 338042
rect 247098 337742 247172 337770
rect 247374 337742 247448 337770
rect 246580 326460 246632 326466
rect 246580 326402 246632 326408
rect 247040 326324 247092 326330
rect 247040 326266 247092 326272
rect 246316 316006 246436 316034
rect 246316 7002 246344 316006
rect 246304 6996 246356 7002
rect 246304 6938 246356 6944
rect 245936 4140 245988 4146
rect 245936 4082 245988 4088
rect 245752 4004 245804 4010
rect 245752 3946 245804 3952
rect 244648 3868 244700 3874
rect 244648 3810 244700 3816
rect 245200 3732 245252 3738
rect 245200 3674 245252 3680
rect 245212 480 245240 3674
rect 247052 3602 247080 326266
rect 247144 6225 247172 337742
rect 247316 326460 247368 326466
rect 247316 326402 247368 326408
rect 247224 326392 247276 326398
rect 247224 326334 247276 326340
rect 247236 6361 247264 326334
rect 247328 10402 247356 326402
rect 247316 10396 247368 10402
rect 247316 10338 247368 10344
rect 247420 10334 247448 337742
rect 247512 326330 247540 338014
rect 247788 326398 247816 338014
rect 248064 326466 248092 338014
rect 248432 336530 248460 338014
rect 248708 336682 248736 338014
rect 248984 336818 249012 338014
rect 248616 336654 248736 336682
rect 248892 336790 249012 336818
rect 248420 336524 248472 336530
rect 248420 336466 248472 336472
rect 248052 326460 248104 326466
rect 248052 326402 248104 326408
rect 247776 326392 247828 326398
rect 247776 326334 247828 326340
rect 248512 326392 248564 326398
rect 248512 326334 248564 326340
rect 247500 326324 247552 326330
rect 247500 326266 247552 326272
rect 248420 12572 248472 12578
rect 248420 12514 248472 12520
rect 248432 10470 248460 12514
rect 248420 10464 248472 10470
rect 248420 10406 248472 10412
rect 247408 10328 247460 10334
rect 247408 10270 247460 10276
rect 247592 6996 247644 7002
rect 247592 6938 247644 6944
rect 247222 6352 247278 6361
rect 247222 6287 247278 6296
rect 247130 6216 247186 6225
rect 247130 6151 247186 6160
rect 247040 3596 247092 3602
rect 247040 3538 247092 3544
rect 246396 3528 246448 3534
rect 246396 3470 246448 3476
rect 246408 480 246436 3470
rect 247604 480 247632 6938
rect 248524 6633 248552 326334
rect 248510 6624 248566 6633
rect 248510 6559 248566 6568
rect 248616 6497 248644 336654
rect 248892 335354 248920 336790
rect 249260 336682 249288 338014
rect 248708 335326 248920 335354
rect 248984 336654 249288 336682
rect 248708 12578 248736 335326
rect 248984 316034 249012 336654
rect 249064 336048 249116 336054
rect 249064 335990 249116 335996
rect 248800 316006 249012 316034
rect 248696 12572 248748 12578
rect 248696 12514 248748 12520
rect 248800 11778 248828 316006
rect 248708 11750 248828 11778
rect 248602 6488 248658 6497
rect 248602 6423 248658 6432
rect 248708 3398 248736 11750
rect 248788 8968 248840 8974
rect 248788 8910 248840 8916
rect 248696 3392 248748 3398
rect 248696 3334 248748 3340
rect 248800 480 248828 8910
rect 249076 4078 249104 335990
rect 249628 326398 249656 338014
rect 249616 326392 249668 326398
rect 249616 326334 249668 326340
rect 249892 326392 249944 326398
rect 249892 326334 249944 326340
rect 249904 10606 249932 326334
rect 249892 10600 249944 10606
rect 249892 10542 249944 10548
rect 249996 10538 250024 338014
rect 250180 336598 250208 338014
rect 250168 336592 250220 336598
rect 250168 336534 250220 336540
rect 250456 316034 250484 338014
rect 250824 326398 250852 338014
rect 251238 337822 251266 338028
rect 251376 338014 251528 338042
rect 251652 338014 251896 338042
rect 252020 338014 252172 338042
rect 252296 338014 252448 338042
rect 252724 338014 252876 338042
rect 251226 337816 251278 337822
rect 251226 337758 251278 337764
rect 250812 326392 250864 326398
rect 250812 326334 250864 326340
rect 251272 326392 251324 326398
rect 251272 326334 251324 326340
rect 250088 316006 250484 316034
rect 249984 10532 250036 10538
rect 249984 10474 250036 10480
rect 250088 6254 250116 316006
rect 251284 7682 251312 326334
rect 251376 7750 251404 338014
rect 251548 337816 251600 337822
rect 251548 337758 251600 337764
rect 251560 328454 251588 337758
rect 251468 328426 251588 328454
rect 251468 321722 251496 328426
rect 251468 321694 251588 321722
rect 251456 320748 251508 320754
rect 251456 320690 251508 320696
rect 251468 10674 251496 320690
rect 251456 10668 251508 10674
rect 251456 10610 251508 10616
rect 251364 7744 251416 7750
rect 251364 7686 251416 7692
rect 251272 7676 251324 7682
rect 251272 7618 251324 7624
rect 251180 7608 251232 7614
rect 251180 7550 251232 7556
rect 250076 6248 250128 6254
rect 250076 6190 250128 6196
rect 249064 4072 249116 4078
rect 249064 4014 249116 4020
rect 249984 3392 250036 3398
rect 249984 3334 250036 3340
rect 249996 480 250024 3334
rect 251192 480 251220 7550
rect 251560 3330 251588 321694
rect 251652 320754 251680 338014
rect 252020 336666 252048 338014
rect 252008 336660 252060 336666
rect 252008 336602 252060 336608
rect 251824 336252 251876 336258
rect 251824 336194 251876 336200
rect 251640 320748 251692 320754
rect 251640 320690 251692 320696
rect 251836 3670 251864 336194
rect 252296 326398 252324 338014
rect 252468 336116 252520 336122
rect 252468 336058 252520 336064
rect 252284 326392 252336 326398
rect 252284 326334 252336 326340
rect 252480 6914 252508 336058
rect 252744 326460 252796 326466
rect 252744 326402 252796 326408
rect 252652 326392 252704 326398
rect 252652 326334 252704 326340
rect 252664 7818 252692 326334
rect 252756 10810 252784 326402
rect 252744 10804 252796 10810
rect 252744 10746 252796 10752
rect 252848 10742 252876 338014
rect 252940 338014 253092 338042
rect 253216 338014 253368 338042
rect 253492 338014 253644 338042
rect 253768 338014 253920 338042
rect 254044 338014 254288 338042
rect 254412 338014 254564 338042
rect 254688 338014 254840 338042
rect 254964 338014 255116 338042
rect 252836 10736 252888 10742
rect 252836 10678 252888 10684
rect 252652 7812 252704 7818
rect 252652 7754 252704 7760
rect 252388 6886 252508 6914
rect 251824 3664 251876 3670
rect 251824 3606 251876 3612
rect 251548 3324 251600 3330
rect 251548 3266 251600 3272
rect 252388 480 252416 6886
rect 252940 3262 252968 338014
rect 253216 326398 253244 338014
rect 253492 326466 253520 338014
rect 253768 336734 253796 338014
rect 253756 336728 253808 336734
rect 253756 336670 253808 336676
rect 253480 326460 253532 326466
rect 253480 326402 253532 326408
rect 253204 326392 253256 326398
rect 253204 326334 253256 326340
rect 254044 6934 254072 338014
rect 254412 335354 254440 338014
rect 254688 336682 254716 338014
rect 254228 335326 254440 335354
rect 254504 336654 254716 336682
rect 254124 330540 254176 330546
rect 254124 330482 254176 330488
rect 254136 12073 254164 330482
rect 254122 12064 254178 12073
rect 254122 11999 254178 12008
rect 254228 11801 254256 335326
rect 254504 316034 254532 336654
rect 254584 336456 254636 336462
rect 254584 336398 254636 336404
rect 254320 316006 254532 316034
rect 254214 11792 254270 11801
rect 254214 11727 254270 11736
rect 254032 6928 254084 6934
rect 254032 6870 254084 6876
rect 253480 3664 253532 3670
rect 253480 3606 253532 3612
rect 252928 3256 252980 3262
rect 252928 3198 252980 3204
rect 253492 480 253520 3606
rect 254320 3194 254348 316006
rect 254596 3738 254624 336398
rect 254964 330546 254992 338014
rect 255470 337770 255498 338028
rect 255608 338014 255760 338042
rect 255884 338014 256036 338042
rect 256160 338014 256312 338042
rect 256436 338014 256680 338042
rect 256804 338014 256956 338042
rect 257080 338014 257232 338042
rect 257356 338014 257508 338042
rect 257632 338014 257876 338042
rect 258152 338014 258304 338042
rect 255470 337742 255544 337770
rect 254952 330540 255004 330546
rect 254952 330482 255004 330488
rect 255412 327684 255464 327690
rect 255412 327626 255464 327632
rect 255424 11762 255452 327626
rect 255516 11937 255544 337742
rect 255608 335986 255636 338014
rect 255596 335980 255648 335986
rect 255596 335922 255648 335928
rect 255884 316034 255912 338014
rect 256160 327690 256188 338014
rect 256436 335850 256464 338014
rect 256608 336388 256660 336394
rect 256608 336330 256660 336336
rect 256424 335844 256476 335850
rect 256424 335786 256476 335792
rect 256148 327684 256200 327690
rect 256148 327626 256200 327632
rect 255608 316006 255912 316034
rect 255502 11928 255558 11937
rect 255502 11863 255558 11872
rect 255412 11756 255464 11762
rect 255412 11698 255464 11704
rect 255608 10878 255636 316006
rect 255596 10872 255648 10878
rect 255596 10814 255648 10820
rect 254676 7676 254728 7682
rect 254676 7618 254728 7624
rect 254584 3732 254636 3738
rect 254584 3674 254636 3680
rect 254308 3188 254360 3194
rect 254308 3130 254360 3136
rect 254688 480 254716 7618
rect 256620 3602 256648 336330
rect 256700 330540 256752 330546
rect 256700 330482 256752 330488
rect 255872 3596 255924 3602
rect 255872 3538 255924 3544
rect 256608 3596 256660 3602
rect 256608 3538 256660 3544
rect 255884 480 255912 3538
rect 256712 3126 256740 330482
rect 256804 10946 256832 338014
rect 256884 326800 256936 326806
rect 256884 326742 256936 326748
rect 256896 11014 256924 326742
rect 257080 316034 257108 338014
rect 257356 330546 257384 338014
rect 257344 330540 257396 330546
rect 257344 330482 257396 330488
rect 257632 326806 257660 338014
rect 258172 336728 258224 336734
rect 258172 336670 258224 336676
rect 257620 326800 257672 326806
rect 257620 326742 257672 326748
rect 256988 316006 257108 316034
rect 256988 11830 257016 316006
rect 256976 11824 257028 11830
rect 256976 11766 257028 11772
rect 256884 11008 256936 11014
rect 256884 10950 256936 10956
rect 256792 10940 256844 10946
rect 256792 10882 256844 10888
rect 258184 10266 258212 336670
rect 258276 11898 258304 338014
rect 258368 338014 258428 338042
rect 258552 338014 258704 338042
rect 258828 338014 259072 338042
rect 259196 338014 259348 338042
rect 259564 338014 259624 338042
rect 259748 338014 259900 338042
rect 260024 338014 260268 338042
rect 260392 338014 260544 338042
rect 260668 338014 260820 338042
rect 258368 335918 258396 338014
rect 258552 336734 258580 338014
rect 258540 336728 258592 336734
rect 258540 336670 258592 336676
rect 258356 335912 258408 335918
rect 258356 335854 258408 335860
rect 258828 335354 258856 338014
rect 258368 335326 258856 335354
rect 258368 11966 258396 335326
rect 259196 316034 259224 338014
rect 258460 316006 259224 316034
rect 258356 11960 258408 11966
rect 258356 11902 258408 11908
rect 258264 11892 258316 11898
rect 258264 11834 258316 11840
rect 258172 10260 258224 10266
rect 258172 10202 258224 10208
rect 258264 7744 258316 7750
rect 258264 7686 258316 7692
rect 257068 3732 257120 3738
rect 257068 3674 257120 3680
rect 256700 3120 256752 3126
rect 256700 3062 256752 3068
rect 257080 480 257108 3674
rect 258276 480 258304 7686
rect 258460 3058 258488 316006
rect 259564 10198 259592 338014
rect 259748 335354 259776 338014
rect 260024 335782 260052 338014
rect 260012 335776 260064 335782
rect 260012 335718 260064 335724
rect 259656 335326 259776 335354
rect 259656 13122 259684 335326
rect 259736 330540 259788 330546
rect 259736 330482 259788 330488
rect 259748 13190 259776 330482
rect 260392 316034 260420 338014
rect 260668 330546 260696 338014
rect 261082 337770 261110 338028
rect 261220 338014 261464 338042
rect 261588 338014 261740 338042
rect 261864 338014 262016 338042
rect 261082 337742 261156 337770
rect 260748 335980 260800 335986
rect 260748 335922 260800 335928
rect 260656 330540 260708 330546
rect 260656 330482 260708 330488
rect 259840 316006 260420 316034
rect 259736 13184 259788 13190
rect 259736 13126 259788 13132
rect 259644 13116 259696 13122
rect 259644 13058 259696 13064
rect 259552 10192 259604 10198
rect 259552 10134 259604 10140
rect 259840 10130 259868 316006
rect 259828 10124 259880 10130
rect 259828 10066 259880 10072
rect 260654 3632 260710 3641
rect 260654 3567 260710 3576
rect 259460 3392 259512 3398
rect 259460 3334 259512 3340
rect 258448 3052 258500 3058
rect 258448 2994 258500 3000
rect 259472 480 259500 3334
rect 260668 480 260696 3567
rect 260760 3398 260788 335922
rect 261128 330818 261156 337742
rect 261116 330812 261168 330818
rect 261116 330754 261168 330760
rect 261220 330698 261248 338014
rect 260944 330670 261248 330698
rect 260944 10062 260972 330670
rect 261116 330608 261168 330614
rect 261116 330550 261168 330556
rect 261024 330540 261076 330546
rect 261024 330482 261076 330488
rect 261036 13258 261064 330482
rect 261024 13252 261076 13258
rect 261024 13194 261076 13200
rect 260932 10056 260984 10062
rect 260932 9998 260984 10004
rect 260748 3392 260800 3398
rect 260748 3334 260800 3340
rect 261128 2990 261156 330550
rect 261588 330546 261616 338014
rect 261864 335714 261892 338014
rect 262278 337770 262306 338028
rect 262600 338014 262660 338042
rect 262784 338014 262936 338042
rect 263060 338014 263212 338042
rect 263336 338014 263488 338042
rect 263612 338014 263856 338042
rect 263980 338014 264132 338042
rect 264256 338014 264408 338042
rect 264532 338014 264684 338042
rect 262278 337742 262352 337770
rect 261852 335708 261904 335714
rect 261852 335650 261904 335656
rect 261576 330540 261628 330546
rect 261576 330482 261628 330488
rect 262324 9994 262352 337742
rect 262496 330540 262548 330546
rect 262496 330482 262548 330488
rect 262404 326596 262456 326602
rect 262404 326538 262456 326544
rect 262312 9988 262364 9994
rect 262312 9930 262364 9936
rect 262416 9926 262444 326538
rect 262508 13394 262536 330482
rect 262496 13388 262548 13394
rect 262496 13330 262548 13336
rect 262600 13326 262628 338014
rect 262784 316034 262812 338014
rect 263060 326602 263088 338014
rect 263336 330546 263364 338014
rect 263508 336592 263560 336598
rect 263508 336534 263560 336540
rect 263324 330540 263376 330546
rect 263324 330482 263376 330488
rect 263048 326596 263100 326602
rect 263048 326538 263100 326544
rect 262692 316006 262812 316034
rect 262588 13320 262640 13326
rect 262588 13262 262640 13268
rect 262404 9920 262456 9926
rect 262404 9862 262456 9868
rect 261760 7812 261812 7818
rect 261760 7754 261812 7760
rect 261116 2984 261168 2990
rect 261116 2926 261168 2932
rect 261772 480 261800 7754
rect 262692 2922 262720 316006
rect 263520 2922 263548 336534
rect 263612 335646 263640 338014
rect 263980 336682 264008 338014
rect 263704 336654 264008 336682
rect 263600 335640 263652 335646
rect 263600 335582 263652 335588
rect 263704 9858 263732 336654
rect 264256 335354 264284 338014
rect 263796 335326 264284 335354
rect 263796 13462 263824 335326
rect 264532 316034 264560 338014
rect 265038 337822 265066 338028
rect 265176 338014 265328 338042
rect 265452 338014 265604 338042
rect 265728 338014 265880 338042
rect 266004 338014 266248 338042
rect 266372 338014 266524 338042
rect 266648 338014 266800 338042
rect 266924 338014 267076 338042
rect 267200 338014 267444 338042
rect 267568 338014 267720 338042
rect 267844 338014 267996 338042
rect 268120 338014 268272 338042
rect 268396 338014 268640 338042
rect 268764 338014 268916 338042
rect 269192 338014 269344 338042
rect 265026 337816 265078 337822
rect 265026 337758 265078 337764
rect 265072 330540 265124 330546
rect 265072 330482 265124 330488
rect 263888 316006 264560 316034
rect 263784 13456 263836 13462
rect 263784 13398 263836 13404
rect 263692 9852 263744 9858
rect 263692 9794 263744 9800
rect 262680 2916 262732 2922
rect 262680 2858 262732 2864
rect 262956 2916 263008 2922
rect 262956 2858 263008 2864
rect 263508 2916 263560 2922
rect 263508 2858 263560 2864
rect 262968 480 262996 2858
rect 263888 2854 263916 316006
rect 265084 9722 265112 330482
rect 265176 13530 265204 338014
rect 265256 337816 265308 337822
rect 265256 337758 265308 337764
rect 265164 13524 265216 13530
rect 265164 13466 265216 13472
rect 265268 9790 265296 337758
rect 265452 335578 265480 338014
rect 265440 335572 265492 335578
rect 265440 335514 265492 335520
rect 265728 330546 265756 338014
rect 266004 335442 266032 338014
rect 266372 335510 266400 338014
rect 266360 335504 266412 335510
rect 266360 335446 266412 335452
rect 265992 335436 266044 335442
rect 265992 335378 266044 335384
rect 265716 330540 265768 330546
rect 265716 330482 265768 330488
rect 266452 330540 266504 330546
rect 266452 330482 266504 330488
rect 265256 9784 265308 9790
rect 265256 9726 265308 9732
rect 265072 9716 265124 9722
rect 265072 9658 265124 9664
rect 266464 6322 266492 330482
rect 266544 330472 266596 330478
rect 266544 330414 266596 330420
rect 266556 7886 266584 330414
rect 266648 12034 266676 338014
rect 266924 330546 266952 338014
rect 266912 330540 266964 330546
rect 266912 330482 266964 330488
rect 267200 330478 267228 338014
rect 267188 330472 267240 330478
rect 267188 330414 267240 330420
rect 267568 316034 267596 338014
rect 267648 336660 267700 336666
rect 267648 336602 267700 336608
rect 266740 316006 267596 316034
rect 266636 12028 266688 12034
rect 266636 11970 266688 11976
rect 266544 7880 266596 7886
rect 266544 7822 266596 7828
rect 266452 6316 266504 6322
rect 266452 6258 266504 6264
rect 266740 4865 266768 316006
rect 266726 4856 266782 4865
rect 266726 4791 266782 4800
rect 265348 3936 265400 3942
rect 265348 3878 265400 3884
rect 264152 3800 264204 3806
rect 264152 3742 264204 3748
rect 263876 2848 263928 2854
rect 263876 2790 263928 2796
rect 264164 480 264192 3742
rect 265360 480 265388 3878
rect 267660 3194 267688 336602
rect 267740 330472 267792 330478
rect 267740 330414 267792 330420
rect 267752 5001 267780 330414
rect 267844 6390 267872 338014
rect 267924 330540 267976 330546
rect 267924 330482 267976 330488
rect 267936 7954 267964 330482
rect 268120 316034 268148 338014
rect 268396 330478 268424 338014
rect 268764 330546 268792 338014
rect 269028 335980 269080 335986
rect 269028 335922 269080 335928
rect 268752 330540 268804 330546
rect 268752 330482 268804 330488
rect 268384 330472 268436 330478
rect 268384 330414 268436 330420
rect 268028 316006 268148 316034
rect 268028 9217 268056 316006
rect 268014 9208 268070 9217
rect 268014 9143 268070 9152
rect 267924 7948 267976 7954
rect 267924 7890 267976 7896
rect 269040 6914 269068 335922
rect 269120 330540 269172 330546
rect 269120 330482 269172 330488
rect 269132 8022 269160 330482
rect 269212 330472 269264 330478
rect 269212 330414 269264 330420
rect 269224 9042 269252 330414
rect 269316 9353 269344 338014
rect 269408 338014 269468 338042
rect 269592 338014 269836 338042
rect 269960 338014 270112 338042
rect 270236 338014 270388 338042
rect 270512 338014 270664 338042
rect 270788 338014 271032 338042
rect 271156 338014 271308 338042
rect 271432 338014 271584 338042
rect 271708 338014 271860 338042
rect 272168 338014 272228 338042
rect 272352 338014 272504 338042
rect 272628 338014 272780 338042
rect 272904 338014 273056 338042
rect 273364 338014 273424 338042
rect 273548 338014 273700 338042
rect 273824 338014 273976 338042
rect 274100 338014 274252 338042
rect 274376 338014 274620 338042
rect 274744 338014 274896 338042
rect 275020 338014 275172 338042
rect 275296 338014 275448 338042
rect 275572 338014 275816 338042
rect 276032 338014 276092 338042
rect 276308 338014 276368 338042
rect 276492 338014 276644 338042
rect 276768 338014 277012 338042
rect 277136 338014 277288 338042
rect 277412 338014 277564 338042
rect 277688 338014 277840 338042
rect 277964 338014 278208 338042
rect 278332 338014 278484 338042
rect 278608 338014 278760 338042
rect 278976 338014 279036 338042
rect 279160 338014 279404 338042
rect 279528 338014 279680 338042
rect 279804 338014 279956 338042
rect 280172 338014 280232 338042
rect 280356 338014 280600 338042
rect 280724 338014 280876 338042
rect 281000 338014 281152 338042
rect 281276 338014 281428 338042
rect 269408 12102 269436 338014
rect 269592 330546 269620 338014
rect 269580 330540 269632 330546
rect 269580 330482 269632 330488
rect 269960 330478 269988 338014
rect 269948 330472 270000 330478
rect 269948 330414 270000 330420
rect 270236 316034 270264 338014
rect 269500 316006 270264 316034
rect 269500 12170 269528 316006
rect 269488 12164 269540 12170
rect 269488 12106 269540 12112
rect 269396 12096 269448 12102
rect 269396 12038 269448 12044
rect 269302 9344 269358 9353
rect 269302 9279 269358 9288
rect 269212 9036 269264 9042
rect 269212 8978 269264 8984
rect 270512 8090 270540 338014
rect 270788 335354 270816 338014
rect 271156 335354 271184 338014
rect 271236 335912 271288 335918
rect 271236 335854 271288 335860
rect 270696 335326 270816 335354
rect 271064 335326 271184 335354
rect 270592 330472 270644 330478
rect 270592 330414 270644 330420
rect 270604 8158 270632 330414
rect 270696 9110 270724 335326
rect 270776 330540 270828 330546
rect 270776 330482 270828 330488
rect 270788 9178 270816 330482
rect 271064 316034 271092 335326
rect 271248 316034 271276 335854
rect 271432 330478 271460 338014
rect 271708 330546 271736 338014
rect 272168 330818 272196 338014
rect 272352 335354 272380 338014
rect 272260 335326 272380 335354
rect 272156 330812 272208 330818
rect 272156 330754 272208 330760
rect 272260 330698 272288 335326
rect 271984 330670 272288 330698
rect 271696 330540 271748 330546
rect 271696 330482 271748 330488
rect 271420 330472 271472 330478
rect 271420 330414 271472 330420
rect 271880 330472 271932 330478
rect 271880 330414 271932 330420
rect 270880 316006 271092 316034
rect 271156 316006 271276 316034
rect 270880 12238 270908 316006
rect 270868 12232 270920 12238
rect 270868 12174 270920 12180
rect 270776 9172 270828 9178
rect 270776 9114 270828 9120
rect 270684 9104 270736 9110
rect 270684 9046 270736 9052
rect 270592 8152 270644 8158
rect 270592 8094 270644 8100
rect 270500 8084 270552 8090
rect 270500 8026 270552 8032
rect 269120 8016 269172 8022
rect 269120 7958 269172 7964
rect 268856 6886 269068 6914
rect 267832 6384 267884 6390
rect 267832 6326 267884 6332
rect 267738 4992 267794 5001
rect 267738 4927 267794 4936
rect 267738 3768 267794 3777
rect 267738 3703 267794 3712
rect 266544 3188 266596 3194
rect 266544 3130 266596 3136
rect 267648 3188 267700 3194
rect 267648 3130 267700 3136
rect 266556 480 266584 3130
rect 267752 480 267780 3703
rect 268856 480 268884 6886
rect 271156 3942 271184 316006
rect 271892 6458 271920 330414
rect 271984 8226 272012 330670
rect 272156 330608 272208 330614
rect 272156 330550 272208 330556
rect 272064 330540 272116 330546
rect 272064 330482 272116 330488
rect 272076 9246 272104 330482
rect 272168 12306 272196 330550
rect 272628 330546 272656 338014
rect 272616 330540 272668 330546
rect 272616 330482 272668 330488
rect 272904 330478 272932 338014
rect 272892 330472 272944 330478
rect 272892 330414 272944 330420
rect 273260 323332 273312 323338
rect 273260 323274 273312 323280
rect 272156 12300 272208 12306
rect 272156 12242 272208 12248
rect 272064 9240 272116 9246
rect 272064 9182 272116 9188
rect 271972 8220 272024 8226
rect 271972 8162 272024 8168
rect 273272 6526 273300 323274
rect 273364 8294 273392 338014
rect 273444 326392 273496 326398
rect 273444 326334 273496 326340
rect 273352 8288 273404 8294
rect 273352 8230 273404 8236
rect 273456 7546 273484 326334
rect 273548 9314 273576 338014
rect 273824 323338 273852 338014
rect 274100 326398 274128 338014
rect 274088 326392 274140 326398
rect 274088 326334 274140 326340
rect 273812 323332 273864 323338
rect 273812 323274 273864 323280
rect 274376 316034 274404 338014
rect 274744 336682 274772 338014
rect 274652 336654 274772 336682
rect 274548 335844 274600 335850
rect 274548 335786 274600 335792
rect 273640 316006 274404 316034
rect 273640 9382 273668 316006
rect 273628 9376 273680 9382
rect 273628 9318 273680 9324
rect 273536 9308 273588 9314
rect 273536 9250 273588 9256
rect 273444 7540 273496 7546
rect 273444 7482 273496 7488
rect 273260 6520 273312 6526
rect 273260 6462 273312 6468
rect 271880 6452 271932 6458
rect 271880 6394 271932 6400
rect 271236 4956 271288 4962
rect 271236 4898 271288 4904
rect 271144 3936 271196 3942
rect 271144 3878 271196 3884
rect 270040 3868 270092 3874
rect 270040 3810 270092 3816
rect 270052 480 270080 3810
rect 271248 480 271276 4898
rect 272432 3936 272484 3942
rect 272432 3878 272484 3884
rect 272444 480 272472 3878
rect 274560 3398 274588 335786
rect 274652 6594 274680 336654
rect 275020 336546 275048 338014
rect 274744 336518 275048 336546
rect 274744 7478 274772 336518
rect 275296 335354 275324 338014
rect 274836 335326 275324 335354
rect 274836 12374 274864 335326
rect 275572 316034 275600 338014
rect 274928 316006 275600 316034
rect 274928 12442 274956 316006
rect 274916 12436 274968 12442
rect 274916 12378 274968 12384
rect 274824 12368 274876 12374
rect 274824 12310 274876 12316
rect 274732 7472 274784 7478
rect 274732 7414 274784 7420
rect 276032 6662 276060 338014
rect 276204 326460 276256 326466
rect 276204 326402 276256 326408
rect 276112 326392 276164 326398
rect 276112 326334 276164 326340
rect 276124 6730 276152 326334
rect 276216 7342 276244 326402
rect 276308 7410 276336 338014
rect 276492 316034 276520 338014
rect 276768 326398 276796 338014
rect 277136 326466 277164 338014
rect 277412 335374 277440 338014
rect 277688 336682 277716 338014
rect 277504 336654 277716 336682
rect 277400 335368 277452 335374
rect 277400 335310 277452 335316
rect 277124 326460 277176 326466
rect 277124 326402 277176 326408
rect 276756 326392 276808 326398
rect 276756 326334 276808 326340
rect 276400 316006 276520 316034
rect 276400 11694 276428 316006
rect 276388 11688 276440 11694
rect 276388 11630 276440 11636
rect 276296 7404 276348 7410
rect 276296 7346 276348 7352
rect 276204 7336 276256 7342
rect 276204 7278 276256 7284
rect 277504 6798 277532 336654
rect 277964 335354 277992 338014
rect 278332 336734 278360 338014
rect 278320 336728 278372 336734
rect 278320 336670 278372 336676
rect 277596 335326 277992 335354
rect 277596 7274 277624 335326
rect 278608 316034 278636 338014
rect 278976 328454 279004 338014
rect 279160 335354 279188 338014
rect 278884 328426 279004 328454
rect 279068 335326 279188 335354
rect 278780 326732 278832 326738
rect 278780 326674 278832 326680
rect 277688 316006 278636 316034
rect 277584 7268 277636 7274
rect 277584 7210 277636 7216
rect 277688 6866 277716 316006
rect 277676 6860 277728 6866
rect 277676 6802 277728 6808
rect 277492 6792 277544 6798
rect 277492 6734 277544 6740
rect 276112 6724 276164 6730
rect 276112 6666 276164 6672
rect 276020 6656 276072 6662
rect 276020 6598 276072 6604
rect 274640 6588 274692 6594
rect 274640 6530 274692 6536
rect 278792 5137 278820 326674
rect 278884 326482 278912 328426
rect 279068 326738 279096 335326
rect 279056 326732 279108 326738
rect 279056 326674 279108 326680
rect 278884 326454 279004 326482
rect 278872 326392 278924 326398
rect 278872 326334 278924 326340
rect 278884 6118 278912 326334
rect 278976 11626 279004 326454
rect 279528 326398 279556 338014
rect 279516 326392 279568 326398
rect 279516 326334 279568 326340
rect 279804 316034 279832 338014
rect 279068 316006 279832 316034
rect 278964 11620 279016 11626
rect 278964 11562 279016 11568
rect 279068 11558 279096 316006
rect 279056 11552 279108 11558
rect 279056 11494 279108 11500
rect 278872 6112 278924 6118
rect 278872 6054 278924 6060
rect 278778 5128 278834 5137
rect 278778 5063 278834 5072
rect 280172 5030 280200 338014
rect 280252 326460 280304 326466
rect 280252 326402 280304 326408
rect 280264 5098 280292 326402
rect 280356 6050 280384 338014
rect 280436 326392 280488 326398
rect 280436 326334 280488 326340
rect 280344 6044 280396 6050
rect 280344 5986 280396 5992
rect 280448 5982 280476 326334
rect 280724 316034 280752 338014
rect 281000 326466 281028 338014
rect 280988 326460 281040 326466
rect 280988 326402 281040 326408
rect 281276 326398 281304 338014
rect 281782 337770 281810 338028
rect 281920 338014 282072 338042
rect 282196 338014 282348 338042
rect 282472 338014 282624 338042
rect 282932 338014 282992 338042
rect 283208 338014 283268 338042
rect 283392 338014 283544 338042
rect 283668 338014 283820 338042
rect 283944 338014 284188 338042
rect 284464 338014 284616 338042
rect 281782 337742 281856 337770
rect 281540 336728 281592 336734
rect 281540 336670 281592 336676
rect 281264 326392 281316 326398
rect 281264 326334 281316 326340
rect 280540 316006 280752 316034
rect 280540 11490 280568 316006
rect 280528 11484 280580 11490
rect 280528 11426 280580 11432
rect 280436 5976 280488 5982
rect 280436 5918 280488 5924
rect 281552 5166 281580 336670
rect 281724 326460 281776 326466
rect 281724 326402 281776 326408
rect 281632 326392 281684 326398
rect 281632 326334 281684 326340
rect 281644 5914 281672 326334
rect 281736 9450 281764 326402
rect 281828 11422 281856 337742
rect 281920 336734 281948 338014
rect 281908 336728 281960 336734
rect 281908 336670 281960 336676
rect 282196 326398 282224 338014
rect 282276 336728 282328 336734
rect 282276 336670 282328 336676
rect 282184 326392 282236 326398
rect 282184 326334 282236 326340
rect 282288 316034 282316 336670
rect 282472 326466 282500 338014
rect 282460 326460 282512 326466
rect 282460 326402 282512 326408
rect 282196 316006 282316 316034
rect 281816 11416 281868 11422
rect 281816 11358 281868 11364
rect 281724 9444 281776 9450
rect 281724 9386 281776 9392
rect 281632 5908 281684 5914
rect 281632 5850 281684 5856
rect 281540 5160 281592 5166
rect 281540 5102 281592 5108
rect 280252 5092 280304 5098
rect 280252 5034 280304 5040
rect 280160 5024 280212 5030
rect 280160 4966 280212 4972
rect 274824 4548 274876 4554
rect 274824 4490 274876 4496
rect 273628 3392 273680 3398
rect 273628 3334 273680 3340
rect 274548 3392 274600 3398
rect 274548 3334 274600 3340
rect 273640 480 273668 3334
rect 274836 480 274864 4490
rect 279516 4140 279568 4146
rect 279516 4082 279568 4088
rect 276020 4072 276072 4078
rect 276020 4014 276072 4020
rect 276032 480 276060 4014
rect 277124 4004 277176 4010
rect 277124 3946 277176 3952
rect 277136 480 277164 3946
rect 278320 3460 278372 3466
rect 278320 3402 278372 3408
rect 278332 480 278360 3402
rect 279528 480 279556 4082
rect 282196 3466 282224 316006
rect 282932 5234 282960 338014
rect 283104 326460 283156 326466
rect 283104 326402 283156 326408
rect 283012 326392 283064 326398
rect 283012 326334 283064 326340
rect 283024 5302 283052 326334
rect 283116 5778 283144 326402
rect 283208 5846 283236 338014
rect 283392 316034 283420 338014
rect 283668 326398 283696 338014
rect 283944 326466 283972 338014
rect 284300 336796 284352 336802
rect 284300 336738 284352 336744
rect 283932 326460 283984 326466
rect 283932 326402 283984 326408
rect 283656 326392 283708 326398
rect 283656 326334 283708 326340
rect 283300 316006 283420 316034
rect 283300 9518 283328 316006
rect 283288 9512 283340 9518
rect 283288 9454 283340 9460
rect 283196 5840 283248 5846
rect 283196 5782 283248 5788
rect 283104 5772 283156 5778
rect 283104 5714 283156 5720
rect 284312 5370 284340 336738
rect 284588 335354 284616 338014
rect 284680 338014 284740 338042
rect 284864 338014 285108 338042
rect 285232 338014 285384 338042
rect 285508 338014 285660 338042
rect 285784 338014 285936 338042
rect 286060 338014 286304 338042
rect 286428 338014 286580 338042
rect 286704 338014 286856 338042
rect 284680 336802 284708 338014
rect 284668 336796 284720 336802
rect 284668 336738 284720 336744
rect 284864 335354 284892 338014
rect 284588 335326 284708 335354
rect 284680 328454 284708 335326
rect 284588 328426 284708 328454
rect 284772 335326 284892 335354
rect 284484 326732 284536 326738
rect 284484 326674 284536 326680
rect 284392 326460 284444 326466
rect 284392 326402 284444 326408
rect 284404 5438 284432 326402
rect 284496 5710 284524 326674
rect 284588 326482 284616 328426
rect 284772 326738 284800 335326
rect 284760 326732 284812 326738
rect 284760 326674 284812 326680
rect 284588 326454 284708 326482
rect 284576 326392 284628 326398
rect 284576 326334 284628 326340
rect 284588 9654 284616 326334
rect 284576 9648 284628 9654
rect 284576 9590 284628 9596
rect 284680 9586 284708 326454
rect 285232 326398 285260 338014
rect 285508 326466 285536 338014
rect 285588 335776 285640 335782
rect 285588 335718 285640 335724
rect 285496 326460 285548 326466
rect 285496 326402 285548 326408
rect 285220 326392 285272 326398
rect 285220 326334 285272 326340
rect 284668 9580 284720 9586
rect 284668 9522 284720 9528
rect 284484 5704 284536 5710
rect 284484 5646 284536 5652
rect 284392 5432 284444 5438
rect 284392 5374 284444 5380
rect 284300 5364 284352 5370
rect 284300 5306 284352 5312
rect 283012 5296 283064 5302
rect 283012 5238 283064 5244
rect 282920 5228 282972 5234
rect 282920 5170 282972 5176
rect 285600 3466 285628 335718
rect 285680 323604 285732 323610
rect 285680 323546 285732 323552
rect 285692 5506 285720 323546
rect 285784 5642 285812 338014
rect 286060 335354 286088 338014
rect 285876 335326 286088 335354
rect 285876 8906 285904 335326
rect 286428 323610 286456 338014
rect 286416 323604 286468 323610
rect 286416 323546 286468 323552
rect 286704 316034 286732 338014
rect 287118 337770 287146 338028
rect 287348 338014 287500 338042
rect 287624 338014 287776 338042
rect 287900 338014 288052 338042
rect 288176 338014 288328 338042
rect 287118 337742 287192 337770
rect 286968 335640 287020 335646
rect 286968 335582 287020 335588
rect 285968 316006 286732 316034
rect 285968 11354 285996 316006
rect 285956 11348 286008 11354
rect 285956 11290 286008 11296
rect 285864 8900 285916 8906
rect 285864 8842 285916 8848
rect 285772 5636 285824 5642
rect 285772 5578 285824 5584
rect 285680 5500 285732 5506
rect 285680 5442 285732 5448
rect 282184 3460 282236 3466
rect 282184 3402 282236 3408
rect 284300 3460 284352 3466
rect 284300 3402 284352 3408
rect 285588 3460 285640 3466
rect 285588 3402 285640 3408
rect 283104 3324 283156 3330
rect 283104 3266 283156 3272
rect 281908 3256 281960 3262
rect 281908 3198 281960 3204
rect 280712 3120 280764 3126
rect 280712 3062 280764 3068
rect 280724 480 280752 3062
rect 281920 480 281948 3198
rect 283116 480 283144 3266
rect 284312 480 284340 3402
rect 285404 3188 285456 3194
rect 285404 3130 285456 3136
rect 285416 480 285444 3130
rect 286612 598 286824 626
rect 286612 480 286640 598
rect 286796 490 286824 598
rect 286980 490 287008 335582
rect 287164 331214 287192 337742
rect 287164 331186 287284 331214
rect 287060 326528 287112 326534
rect 287060 326470 287112 326476
rect 287072 4758 287100 326470
rect 287152 321836 287204 321842
rect 287152 321778 287204 321784
rect 287060 4752 287112 4758
rect 287060 4694 287112 4700
rect 287164 4690 287192 321778
rect 287256 8838 287284 331186
rect 287348 326534 287376 338014
rect 287336 326528 287388 326534
rect 287336 326470 287388 326476
rect 287336 326392 287388 326398
rect 287336 326334 287388 326340
rect 287244 8832 287296 8838
rect 287244 8774 287296 8780
rect 287348 8770 287376 326334
rect 287624 316034 287652 338014
rect 287900 326398 287928 338014
rect 287888 326392 287940 326398
rect 287888 326334 287940 326340
rect 288176 321842 288204 338014
rect 288682 337770 288710 338028
rect 288820 338014 288972 338042
rect 289096 338014 289248 338042
rect 289372 338014 289524 338042
rect 289892 338014 290044 338042
rect 288682 337742 288756 337770
rect 288348 335708 288400 335714
rect 288348 335650 288400 335656
rect 288164 321836 288216 321842
rect 288164 321778 288216 321784
rect 287440 316006 287652 316034
rect 287440 11286 287468 316006
rect 287428 11280 287480 11286
rect 287428 11222 287480 11228
rect 287336 8764 287388 8770
rect 287336 8706 287388 8712
rect 287152 4684 287204 4690
rect 287152 4626 287204 4632
rect 288360 3466 288388 335650
rect 288728 326874 288756 337742
rect 288716 326868 288768 326874
rect 288716 326810 288768 326816
rect 288716 326664 288768 326670
rect 288716 326606 288768 326612
rect 288440 326460 288492 326466
rect 288440 326402 288492 326408
rect 288452 4622 288480 326402
rect 288624 326392 288676 326398
rect 288624 326334 288676 326340
rect 288532 323604 288584 323610
rect 288532 323546 288584 323552
rect 288544 8702 288572 323546
rect 288636 11150 288664 326334
rect 288728 11218 288756 326606
rect 288820 323610 288848 338014
rect 289096 326466 289124 338014
rect 289084 326460 289136 326466
rect 289084 326402 289136 326408
rect 289372 326398 289400 338014
rect 289728 335572 289780 335578
rect 289728 335514 289780 335520
rect 289360 326392 289412 326398
rect 289360 326334 289412 326340
rect 288808 323604 288860 323610
rect 288808 323546 288860 323552
rect 288716 11212 288768 11218
rect 288716 11154 288768 11160
rect 288624 11144 288676 11150
rect 288624 11086 288676 11092
rect 288532 8696 288584 8702
rect 288532 8638 288584 8644
rect 288440 4616 288492 4622
rect 288440 4558 288492 4564
rect 289740 3466 289768 335514
rect 289912 326392 289964 326398
rect 289912 326334 289964 326340
rect 289924 8566 289952 326334
rect 290016 8634 290044 338014
rect 290108 338014 290168 338042
rect 290292 338014 290444 338042
rect 290568 338014 290720 338042
rect 290844 338014 291088 338042
rect 290108 336190 290136 338014
rect 290292 336326 290320 338014
rect 290280 336320 290332 336326
rect 290280 336262 290332 336268
rect 290096 336184 290148 336190
rect 290096 336126 290148 336132
rect 290568 326398 290596 338014
rect 290556 326392 290608 326398
rect 290556 326334 290608 326340
rect 290844 316034 290872 338014
rect 291350 337770 291378 338028
rect 291580 338014 291640 338042
rect 291764 338014 291916 338042
rect 292040 338014 292284 338042
rect 292408 338014 292560 338042
rect 292684 338014 292836 338042
rect 292960 338014 293112 338042
rect 293236 338014 293480 338042
rect 293604 338014 293756 338042
rect 291350 337742 291424 337770
rect 291200 326460 291252 326466
rect 291200 326402 291252 326408
rect 290108 316006 290872 316034
rect 290004 8628 290056 8634
rect 290004 8570 290056 8576
rect 289912 8560 289964 8566
rect 289912 8502 289964 8508
rect 290108 4486 290136 316006
rect 290096 4480 290148 4486
rect 290096 4422 290148 4428
rect 291212 4418 291240 326402
rect 291292 326324 291344 326330
rect 291292 326266 291344 326272
rect 291304 5574 291332 326266
rect 291396 7206 291424 337742
rect 291476 326392 291528 326398
rect 291476 326334 291528 326340
rect 291488 8430 291516 326334
rect 291580 8498 291608 338014
rect 291764 326466 291792 338014
rect 291752 326460 291804 326466
rect 291752 326402 291804 326408
rect 292040 326330 292068 338014
rect 292408 326398 292436 338014
rect 292396 326392 292448 326398
rect 292396 326334 292448 326340
rect 292028 326324 292080 326330
rect 292028 326266 292080 326272
rect 292580 324284 292632 324290
rect 292580 324226 292632 324232
rect 291568 8492 291620 8498
rect 291568 8434 291620 8440
rect 291476 8424 291528 8430
rect 291476 8366 291528 8372
rect 291384 7200 291436 7206
rect 291384 7142 291436 7148
rect 291292 5568 291344 5574
rect 291292 5510 291344 5516
rect 291200 4412 291252 4418
rect 291200 4354 291252 4360
rect 292592 4282 292620 324226
rect 292684 4350 292712 338014
rect 292960 335354 292988 338014
rect 292776 335326 292988 335354
rect 292776 7138 292804 335326
rect 293236 316034 293264 338014
rect 293604 324290 293632 338014
rect 294018 337770 294046 338028
rect 294156 338014 294308 338042
rect 294432 338014 294676 338042
rect 294800 338014 294952 338042
rect 295076 338014 295228 338042
rect 294018 337742 294092 337770
rect 293960 336796 294012 336802
rect 293960 336738 294012 336744
rect 293868 326732 293920 326738
rect 293868 326674 293920 326680
rect 293880 326210 293908 326674
rect 293972 326380 294000 336738
rect 294064 326534 294092 337742
rect 294052 326528 294104 326534
rect 294052 326470 294104 326476
rect 293972 326352 294092 326380
rect 293880 326182 294000 326210
rect 293592 324284 293644 324290
rect 293592 324226 293644 324232
rect 292868 316006 293264 316034
rect 292868 8362 292896 316006
rect 292856 8356 292908 8362
rect 292856 8298 292908 8304
rect 292764 7132 292816 7138
rect 292764 7074 292816 7080
rect 292672 4344 292724 4350
rect 292672 4286 292724 4292
rect 292580 4276 292632 4282
rect 292580 4218 292632 4224
rect 293972 4214 294000 326182
rect 294064 4894 294092 326352
rect 294052 4888 294104 4894
rect 294052 4830 294104 4836
rect 294156 4826 294184 338014
rect 294432 326738 294460 338014
rect 294800 336802 294828 338014
rect 294788 336796 294840 336802
rect 294788 336738 294840 336744
rect 295076 335354 295104 338014
rect 295490 337770 295518 338028
rect 295628 338014 295872 338042
rect 295996 338014 296148 338042
rect 296272 338014 296424 338042
rect 296548 338014 296700 338042
rect 296824 338014 297068 338042
rect 297192 338014 297344 338042
rect 297468 338014 297620 338042
rect 297744 338014 297896 338042
rect 298204 338014 298264 338042
rect 298388 338014 298540 338042
rect 298664 338014 298816 338042
rect 298940 338014 299092 338042
rect 299216 338014 299460 338042
rect 299584 338014 299736 338042
rect 299860 338014 300012 338042
rect 300136 338014 300288 338042
rect 300412 338014 300656 338042
rect 295490 337742 295564 337770
rect 294524 335326 295104 335354
rect 294420 326732 294472 326738
rect 294420 326674 294472 326680
rect 294524 326618 294552 335326
rect 294248 326590 294552 326618
rect 294248 6186 294276 326590
rect 295536 326534 295564 337742
rect 294328 326528 294380 326534
rect 294328 326470 294380 326476
rect 295524 326528 295576 326534
rect 295524 326470 295576 326476
rect 294340 7070 294368 326470
rect 295628 323762 295656 338014
rect 295996 336258 296024 338014
rect 295984 336252 296036 336258
rect 295984 336194 296036 336200
rect 295444 323734 295656 323762
rect 294328 7064 294380 7070
rect 294328 7006 294380 7012
rect 294236 6180 294288 6186
rect 294236 6122 294288 6128
rect 294144 4820 294196 4826
rect 294144 4762 294196 4768
rect 293960 4208 294012 4214
rect 293960 4150 294012 4156
rect 295444 3505 295472 323734
rect 295524 323604 295576 323610
rect 295524 323546 295576 323552
rect 295430 3496 295486 3505
rect 287796 3460 287848 3466
rect 287796 3402 287848 3408
rect 288348 3460 288400 3466
rect 288348 3402 288400 3408
rect 288992 3460 289044 3466
rect 288992 3402 289044 3408
rect 289728 3460 289780 3466
rect 295430 3431 295486 3440
rect 289728 3402 289780 3408
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 212142 -960 212254 480
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215638 -960 215750 480
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220422 -960 220534 480
rect 221526 -960 221638 480
rect 222722 -960 222834 480
rect 223918 -960 224030 480
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228702 -960 228814 480
rect 229806 -960 229918 480
rect 231002 -960 231114 480
rect 232198 -960 232310 480
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236982 -960 237094 480
rect 238086 -960 238198 480
rect 239282 -960 239394 480
rect 240478 -960 240590 480
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 246366 -960 246478 480
rect 247562 -960 247674 480
rect 248758 -960 248870 480
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254646 -960 254758 480
rect 255842 -960 255954 480
rect 257038 -960 257150 480
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262926 -960 263038 480
rect 264122 -960 264234 480
rect 265318 -960 265430 480
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268814 -960 268926 480
rect 270010 -960 270122 480
rect 271206 -960 271318 480
rect 272402 -960 272514 480
rect 273598 -960 273710 480
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 277094 -960 277206 480
rect 278290 -960 278402 480
rect 279486 -960 279598 480
rect 280682 -960 280794 480
rect 281878 -960 281990 480
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 285374 -960 285486 480
rect 286570 -960 286682 480
rect 286796 462 287008 490
rect 287808 480 287836 3402
rect 289004 480 289032 3402
rect 295536 3369 295564 323546
rect 296272 316034 296300 338014
rect 296548 336054 296576 338014
rect 296824 336462 296852 338014
rect 296812 336456 296864 336462
rect 296812 336398 296864 336404
rect 296536 336048 296588 336054
rect 296536 335990 296588 335996
rect 296904 326460 296956 326466
rect 296904 326402 296956 326408
rect 296812 326392 296864 326398
rect 296812 326334 296864 326340
rect 295720 316006 296300 316034
rect 295720 3466 295748 316006
rect 296824 7002 296852 326334
rect 296916 8974 296944 326402
rect 297192 316034 297220 338014
rect 297468 326398 297496 338014
rect 297744 326466 297772 338014
rect 297732 326460 297784 326466
rect 297732 326402 297784 326408
rect 297456 326392 297508 326398
rect 297456 326334 297508 326340
rect 297008 316006 297220 316034
rect 296904 8968 296956 8974
rect 296904 8910 296956 8916
rect 296812 6996 296864 7002
rect 296812 6938 296864 6944
rect 297008 3534 297036 316006
rect 298204 3602 298232 338014
rect 298284 326392 298336 326398
rect 298284 326334 298336 326340
rect 298296 7682 298324 326334
rect 298284 7676 298336 7682
rect 298284 7618 298336 7624
rect 298388 7614 298416 338014
rect 298664 336122 298692 338014
rect 298652 336116 298704 336122
rect 298652 336058 298704 336064
rect 298940 316034 298968 338014
rect 299216 326398 299244 338014
rect 299584 336394 299612 338014
rect 299572 336388 299624 336394
rect 299572 336330 299624 336336
rect 299204 326392 299256 326398
rect 299204 326334 299256 326340
rect 299572 326392 299624 326398
rect 299572 326334 299624 326340
rect 298480 316006 298968 316034
rect 298376 7608 298428 7614
rect 298376 7550 298428 7556
rect 298480 3670 298508 316006
rect 299584 7750 299612 326334
rect 299860 316034 299888 338014
rect 300136 326398 300164 338014
rect 300412 336530 300440 338014
rect 300918 337770 300946 338028
rect 301056 338014 301208 338042
rect 301332 338014 301484 338042
rect 301608 338014 301852 338042
rect 301976 338014 302128 338042
rect 302252 338014 302404 338042
rect 302528 338014 302680 338042
rect 302804 338014 303048 338042
rect 303172 338014 303324 338042
rect 303448 338014 303600 338042
rect 303724 338014 303876 338042
rect 304000 338014 304244 338042
rect 304368 338014 304520 338042
rect 304644 338014 304796 338042
rect 300918 337742 300992 337770
rect 300400 336524 300452 336530
rect 300400 336466 300452 336472
rect 300124 326392 300176 326398
rect 300124 326334 300176 326340
rect 299676 316006 299888 316034
rect 299572 7744 299624 7750
rect 299572 7686 299624 7692
rect 299676 3738 299704 316006
rect 299664 3732 299716 3738
rect 299664 3674 299716 3680
rect 298468 3664 298520 3670
rect 298468 3606 298520 3612
rect 298560 3664 298612 3670
rect 300964 3641 300992 337742
rect 301056 7818 301084 338014
rect 301332 336598 301360 338014
rect 301320 336592 301372 336598
rect 301320 336534 301372 336540
rect 301608 316034 301636 338014
rect 301976 335918 302004 338014
rect 302252 336666 302280 338014
rect 302240 336660 302292 336666
rect 302240 336602 302292 336608
rect 301964 335912 302016 335918
rect 301964 335854 302016 335860
rect 302424 330540 302476 330546
rect 302424 330482 302476 330488
rect 302332 328976 302384 328982
rect 302332 328918 302384 328924
rect 301148 316006 301636 316034
rect 301044 7812 301096 7818
rect 301044 7754 301096 7760
rect 301148 3806 301176 316006
rect 302344 3874 302372 328918
rect 302436 4962 302464 330482
rect 302424 4956 302476 4962
rect 302424 4898 302476 4904
rect 302332 3868 302384 3874
rect 302332 3810 302384 3816
rect 301136 3800 301188 3806
rect 301136 3742 301188 3748
rect 301964 3800 302016 3806
rect 302528 3777 302556 338014
rect 302804 335986 302832 338014
rect 302792 335980 302844 335986
rect 302792 335922 302844 335928
rect 303172 328982 303200 338014
rect 303448 330546 303476 338014
rect 303528 336048 303580 336054
rect 303528 335990 303580 335996
rect 303436 330540 303488 330546
rect 303436 330482 303488 330488
rect 303160 328976 303212 328982
rect 303160 328918 303212 328924
rect 301964 3742 302016 3748
rect 302514 3768 302570 3777
rect 298560 3606 298612 3612
rect 300950 3632 301006 3641
rect 298192 3596 298244 3602
rect 298192 3538 298244 3544
rect 296996 3528 297048 3534
rect 296996 3470 297048 3476
rect 297272 3528 297324 3534
rect 297272 3470 297324 3476
rect 295708 3460 295760 3466
rect 295708 3402 295760 3408
rect 296076 3460 296128 3466
rect 296076 3402 296128 3408
rect 295522 3360 295578 3369
rect 295522 3295 295578 3304
rect 290188 3052 290240 3058
rect 290188 2994 290240 3000
rect 293684 3052 293736 3058
rect 293684 2994 293736 3000
rect 290200 480 290228 2994
rect 291384 2984 291436 2990
rect 291384 2926 291436 2932
rect 291396 480 291424 2926
rect 292580 2848 292632 2854
rect 292580 2790 292632 2796
rect 292592 480 292620 2790
rect 293696 480 293724 2994
rect 294880 2916 294932 2922
rect 294880 2858 294932 2864
rect 294892 480 294920 2858
rect 296088 480 296116 3402
rect 297284 480 297312 3470
rect 298572 1850 298600 3606
rect 300768 3596 300820 3602
rect 300950 3567 301006 3576
rect 300768 3538 300820 3544
rect 299664 3392 299716 3398
rect 299664 3334 299716 3340
rect 298480 1822 298600 1850
rect 298480 480 298508 1822
rect 299676 480 299704 3334
rect 300780 480 300808 3538
rect 301976 480 302004 3742
rect 302514 3703 302570 3712
rect 303172 598 303384 626
rect 303172 480 303200 598
rect 303356 490 303384 598
rect 303540 490 303568 335990
rect 303724 3942 303752 338014
rect 304000 335850 304028 338014
rect 303988 335844 304040 335850
rect 303988 335786 304040 335792
rect 304368 335354 304396 338014
rect 303816 335326 304396 335354
rect 303816 4554 303844 335326
rect 304644 316034 304672 338014
rect 305058 337770 305086 338028
rect 305196 338014 305440 338042
rect 305564 338014 305716 338042
rect 305840 338014 305992 338042
rect 306116 338014 306268 338042
rect 306484 338014 306636 338042
rect 306760 338014 306912 338042
rect 307036 338014 307188 338042
rect 307312 338014 307464 338042
rect 307772 338014 307832 338042
rect 307956 338014 308108 338042
rect 308232 338014 308384 338042
rect 308508 338014 308660 338042
rect 308784 338014 309028 338042
rect 309304 338014 309456 338042
rect 305058 337742 305132 337770
rect 303908 316006 304672 316034
rect 303804 4548 303856 4554
rect 303804 4490 303856 4496
rect 303908 4078 303936 316006
rect 303896 4072 303948 4078
rect 303896 4014 303948 4020
rect 305104 4010 305132 337742
rect 305196 336734 305224 338014
rect 305184 336728 305236 336734
rect 305184 336670 305236 336676
rect 305564 335354 305592 338014
rect 305380 335326 305592 335354
rect 305184 330540 305236 330546
rect 305184 330482 305236 330488
rect 305092 4004 305144 4010
rect 305092 3946 305144 3952
rect 303712 3936 303764 3942
rect 303712 3878 303764 3884
rect 304356 3868 304408 3874
rect 304356 3810 304408 3816
rect 287766 -960 287878 480
rect 288962 -960 289074 480
rect 290158 -960 290270 480
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293654 -960 293766 480
rect 294850 -960 294962 480
rect 296046 -960 296158 480
rect 297242 -960 297354 480
rect 298438 -960 298550 480
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301934 -960 302046 480
rect 303130 -960 303242 480
rect 303356 462 303568 490
rect 304368 480 304396 3810
rect 305196 3194 305224 330482
rect 305380 316034 305408 335326
rect 305840 330546 305868 338014
rect 305828 330540 305880 330546
rect 305828 330482 305880 330488
rect 306116 316034 306144 338014
rect 305288 316006 305408 316034
rect 305472 316006 306144 316034
rect 305288 4146 305316 316006
rect 305276 4140 305328 4146
rect 305276 4082 305328 4088
rect 305472 3738 305500 316006
rect 305552 3936 305604 3942
rect 305552 3878 305604 3884
rect 305460 3732 305512 3738
rect 305460 3674 305512 3680
rect 305184 3188 305236 3194
rect 305184 3130 305236 3136
rect 305564 480 305592 3878
rect 306484 3194 306512 338014
rect 306760 335782 306788 338014
rect 306748 335776 306800 335782
rect 306748 335718 306800 335724
rect 307036 316034 307064 338014
rect 307312 335646 307340 338014
rect 307668 336524 307720 336530
rect 307668 336466 307720 336472
rect 307300 335640 307352 335646
rect 307300 335582 307352 335588
rect 306576 316006 307064 316034
rect 306472 3188 306524 3194
rect 306472 3130 306524 3136
rect 306576 3126 306604 316006
rect 307680 3534 307708 336466
rect 307772 335714 307800 338014
rect 307760 335708 307812 335714
rect 307760 335650 307812 335656
rect 307956 335578 307984 338014
rect 307944 335572 307996 335578
rect 307944 335514 307996 335520
rect 307852 330540 307904 330546
rect 307852 330482 307904 330488
rect 306748 3528 306800 3534
rect 306748 3470 306800 3476
rect 307668 3528 307720 3534
rect 307668 3470 307720 3476
rect 306564 3120 306616 3126
rect 306564 3062 306616 3068
rect 306760 480 306788 3470
rect 307864 2990 307892 330482
rect 307944 330472 307996 330478
rect 307944 330414 307996 330420
rect 307956 4146 307984 330414
rect 307944 4140 307996 4146
rect 307944 4082 307996 4088
rect 307944 3392 307996 3398
rect 307944 3334 307996 3340
rect 307852 2984 307904 2990
rect 307852 2926 307904 2932
rect 307956 480 307984 3334
rect 308232 2854 308260 338014
rect 308508 330546 308536 338014
rect 308496 330540 308548 330546
rect 308496 330482 308548 330488
rect 308784 330478 308812 338014
rect 309140 330608 309192 330614
rect 309140 330550 309192 330556
rect 308772 330472 308824 330478
rect 308772 330414 308824 330420
rect 309152 3670 309180 330550
rect 309232 330540 309284 330546
rect 309232 330482 309284 330488
rect 309140 3664 309192 3670
rect 309140 3606 309192 3612
rect 309244 3534 309272 330482
rect 309324 330472 309376 330478
rect 309324 330414 309376 330420
rect 309336 3602 309364 330414
rect 309324 3596 309376 3602
rect 309324 3538 309376 3544
rect 309232 3528 309284 3534
rect 309232 3470 309284 3476
rect 309048 3460 309100 3466
rect 309048 3402 309100 3408
rect 308220 2848 308272 2854
rect 308220 2790 308272 2796
rect 309060 480 309088 3402
rect 309428 3058 309456 338014
rect 309520 338014 309580 338042
rect 309704 338014 309856 338042
rect 309980 338014 310224 338042
rect 310348 338014 310500 338042
rect 310624 338014 310776 338042
rect 310900 338014 311052 338042
rect 311176 338014 311420 338042
rect 311544 338014 311696 338042
rect 311912 338014 311972 338042
rect 312096 338014 312248 338042
rect 312372 338014 312616 338042
rect 312740 338014 312892 338042
rect 313016 338014 313168 338042
rect 309416 3052 309468 3058
rect 309416 2994 309468 3000
rect 309520 2922 309548 338014
rect 309704 330546 309732 338014
rect 309692 330540 309744 330546
rect 309692 330482 309744 330488
rect 309980 330478 310008 338014
rect 310348 330614 310376 338014
rect 310336 330608 310388 330614
rect 310336 330550 310388 330556
rect 309968 330472 310020 330478
rect 309968 330414 310020 330420
rect 310624 3330 310652 338014
rect 310900 335354 310928 338014
rect 311176 336682 311204 338014
rect 310716 335326 310928 335354
rect 311084 336654 311204 336682
rect 310716 3738 310744 335326
rect 311084 316034 311112 336654
rect 311164 336592 311216 336598
rect 311164 336534 311216 336540
rect 310808 316006 311112 316034
rect 310808 3806 310836 316006
rect 311176 3874 311204 336534
rect 311544 336054 311572 338014
rect 311912 336598 311940 338014
rect 312096 336682 312124 338014
rect 312004 336654 312124 336682
rect 311900 336592 311952 336598
rect 311900 336534 311952 336540
rect 311532 336048 311584 336054
rect 311532 335990 311584 335996
rect 312004 3942 312032 336654
rect 312372 336530 312400 338014
rect 312360 336524 312412 336530
rect 312360 336466 312412 336472
rect 312740 335354 312768 338014
rect 312096 335326 312768 335354
rect 311992 3936 312044 3942
rect 311992 3878 312044 3884
rect 311164 3868 311216 3874
rect 311164 3810 311216 3816
rect 310796 3800 310848 3806
rect 310796 3742 310848 3748
rect 310704 3732 310756 3738
rect 310704 3674 310756 3680
rect 312096 3398 312124 335326
rect 313016 316034 313044 338014
rect 313430 337770 313458 338028
rect 313568 338014 313812 338042
rect 313936 338014 314088 338042
rect 314212 338014 314364 338042
rect 314580 338014 314640 338042
rect 315008 338014 315160 338042
rect 315284 338014 315436 338042
rect 315560 338014 315712 338042
rect 315836 338014 315988 338042
rect 313430 337742 313504 337770
rect 313372 336728 313424 336734
rect 313372 336670 313424 336676
rect 313280 330540 313332 330546
rect 313280 330482 313332 330488
rect 312188 316006 313044 316034
rect 312188 3466 312216 316006
rect 313292 3534 313320 330482
rect 313280 3528 313332 3534
rect 313280 3470 313332 3476
rect 312176 3460 312228 3466
rect 312176 3402 312228 3408
rect 312084 3392 312136 3398
rect 312084 3334 312136 3340
rect 313384 3330 313412 336670
rect 310612 3324 310664 3330
rect 310612 3266 310664 3272
rect 311440 3324 311492 3330
rect 311440 3266 311492 3272
rect 313372 3324 313424 3330
rect 313372 3266 313424 3272
rect 310244 3052 310296 3058
rect 310244 2994 310296 3000
rect 309508 2916 309560 2922
rect 309508 2858 309560 2864
rect 310256 480 310284 2994
rect 311452 480 311480 3266
rect 313476 3058 313504 337742
rect 313568 336734 313596 338014
rect 313556 336728 313608 336734
rect 313556 336670 313608 336676
rect 313936 316034 313964 338014
rect 314212 330546 314240 338014
rect 314580 335354 314608 338014
rect 315132 335646 315160 338014
rect 315408 336326 315436 338014
rect 315396 336320 315448 336326
rect 315396 336262 315448 336268
rect 315120 335640 315172 335646
rect 315120 335582 315172 335588
rect 315684 335374 315712 338014
rect 315960 336122 315988 338014
rect 316144 338014 316204 338042
rect 316480 338014 316632 338042
rect 316756 338014 316908 338042
rect 317032 338014 317276 338042
rect 315948 336116 316000 336122
rect 315948 336058 316000 336064
rect 316144 336054 316172 338014
rect 316604 336530 316632 338014
rect 316592 336524 316644 336530
rect 316592 336466 316644 336472
rect 316880 336462 316908 338014
rect 316868 336456 316920 336462
rect 316868 336398 316920 336404
rect 316316 336320 316368 336326
rect 316316 336262 316368 336268
rect 316132 336048 316184 336054
rect 316132 335990 316184 335996
rect 316132 335640 316184 335646
rect 316132 335582 316184 335588
rect 315672 335368 315724 335374
rect 314580 335326 314700 335354
rect 314200 330540 314252 330546
rect 314200 330482 314252 330488
rect 313568 316006 313964 316034
rect 313464 3052 313516 3058
rect 313464 2994 313516 3000
rect 313568 2922 313596 316006
rect 313832 3528 313884 3534
rect 313832 3470 313884 3476
rect 312636 2916 312688 2922
rect 312636 2858 312688 2864
rect 313556 2916 313608 2922
rect 313556 2858 313608 2864
rect 312648 480 312676 2858
rect 313844 480 313872 3470
rect 314672 490 314700 335326
rect 315672 335310 315724 335316
rect 316144 16574 316172 335582
rect 316328 16574 316356 336262
rect 316144 16546 316264 16574
rect 316328 16546 317184 16574
rect 314856 598 315068 626
rect 314856 490 314884 598
rect 304326 -960 304438 480
rect 305522 -960 305634 480
rect 306718 -960 306830 480
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 310214 -960 310326 480
rect 311410 -960 311522 480
rect 312606 -960 312718 480
rect 313802 -960 313914 480
rect 314672 462 314884 490
rect 315040 480 315068 598
rect 316236 480 316264 16546
rect 317156 2802 317184 16546
rect 317248 2922 317276 338014
rect 317340 338014 317400 338042
rect 317676 338014 317828 338042
rect 317952 338014 318104 338042
rect 318228 338014 318472 338042
rect 318596 338014 318748 338042
rect 318872 338014 319024 338042
rect 319148 338014 319300 338042
rect 319424 338014 319668 338042
rect 319792 338014 319944 338042
rect 317340 3602 317368 338014
rect 317800 336734 317828 338014
rect 317788 336728 317840 336734
rect 317788 336670 317840 336676
rect 318076 336598 318104 338014
rect 318444 336682 318472 338014
rect 318720 336818 318748 338014
rect 318720 336790 318840 336818
rect 318444 336654 318748 336682
rect 318812 336666 318840 336790
rect 318064 336592 318116 336598
rect 318064 336534 318116 336540
rect 318616 336592 318668 336598
rect 318616 336534 318668 336540
rect 317972 336048 318024 336054
rect 317972 335990 318024 335996
rect 317512 335368 317564 335374
rect 317512 335310 317564 335316
rect 317524 6914 317552 335310
rect 317984 325694 318012 335990
rect 317984 325666 318104 325694
rect 318076 16574 318104 325666
rect 318076 16546 318196 16574
rect 317524 6886 318104 6914
rect 317328 3596 317380 3602
rect 317328 3538 317380 3544
rect 317236 2916 317288 2922
rect 317236 2858 317288 2864
rect 317156 2774 317368 2802
rect 317340 480 317368 2774
rect 318076 490 318104 6886
rect 318168 3126 318196 16546
rect 318628 3398 318656 336534
rect 318616 3392 318668 3398
rect 318616 3334 318668 3340
rect 318720 3330 318748 336654
rect 318800 336660 318852 336666
rect 318800 336602 318852 336608
rect 318892 336116 318944 336122
rect 318892 336058 318944 336064
rect 318904 16574 318932 336058
rect 318996 335442 319024 338014
rect 319272 336258 319300 338014
rect 319260 336252 319312 336258
rect 319260 336194 319312 336200
rect 319640 335578 319668 338014
rect 319916 336326 319944 338014
rect 320008 338014 320068 338042
rect 320344 338014 320496 338042
rect 320620 338014 320772 338042
rect 320988 338014 321140 338042
rect 320008 336394 320036 338014
rect 319996 336388 320048 336394
rect 319996 336330 320048 336336
rect 319904 336320 319956 336326
rect 319904 336262 319956 336268
rect 319628 335572 319680 335578
rect 319628 335514 319680 335520
rect 320088 335572 320140 335578
rect 320088 335514 320140 335520
rect 318984 335436 319036 335442
rect 318984 335378 319036 335384
rect 318904 16546 319760 16574
rect 318708 3324 318760 3330
rect 318708 3266 318760 3272
rect 318156 3120 318208 3126
rect 318156 3062 318208 3068
rect 318352 598 318564 626
rect 318352 490 318380 598
rect 314998 -960 315110 480
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318076 462 318380 490
rect 318536 480 318564 598
rect 319732 480 319760 16546
rect 320100 4078 320128 335514
rect 320468 330478 320496 338014
rect 320744 336190 320772 338014
rect 320824 336728 320876 336734
rect 320824 336670 320876 336676
rect 320732 336184 320784 336190
rect 320732 336126 320784 336132
rect 320456 330472 320508 330478
rect 320456 330414 320508 330420
rect 320088 4072 320140 4078
rect 320088 4014 320140 4020
rect 320836 3874 320864 336670
rect 320916 336524 320968 336530
rect 320916 336466 320968 336472
rect 320824 3868 320876 3874
rect 320824 3810 320876 3816
rect 320928 3534 320956 336466
rect 321112 336122 321140 338014
rect 321204 338014 321264 338042
rect 321388 338014 321540 338042
rect 321816 338014 322060 338042
rect 322184 338014 322336 338042
rect 322460 338014 322612 338042
rect 322736 338014 322888 338042
rect 323012 338014 323256 338042
rect 323380 338014 323532 338042
rect 323656 338014 323808 338042
rect 321204 336734 321232 338014
rect 321192 336728 321244 336734
rect 321192 336670 321244 336676
rect 321100 336116 321152 336122
rect 321100 336058 321152 336064
rect 321388 330562 321416 338014
rect 322032 336734 322060 338014
rect 321468 336728 321520 336734
rect 321468 336670 321520 336676
rect 322020 336728 322072 336734
rect 322020 336670 322072 336676
rect 321296 330534 321416 330562
rect 321296 3738 321324 330534
rect 321376 330472 321428 330478
rect 321376 330414 321428 330420
rect 321284 3732 321336 3738
rect 321284 3674 321336 3680
rect 321388 3670 321416 330414
rect 321376 3664 321428 3670
rect 321376 3606 321428 3612
rect 320916 3528 320968 3534
rect 320916 3470 320968 3476
rect 320916 3120 320968 3126
rect 320916 3062 320968 3068
rect 320928 480 320956 3062
rect 321480 2990 321508 336670
rect 322204 336660 322256 336666
rect 322204 336602 322256 336608
rect 322216 3806 322244 336602
rect 322308 335510 322336 338014
rect 322388 336456 322440 336462
rect 322388 336398 322440 336404
rect 322296 335504 322348 335510
rect 322296 335446 322348 335452
rect 322400 316034 322428 336398
rect 322584 335354 322612 338014
rect 322756 336728 322808 336734
rect 322756 336670 322808 336676
rect 322584 335326 322704 335354
rect 322308 316006 322428 316034
rect 322204 3800 322256 3806
rect 322204 3742 322256 3748
rect 322308 3534 322336 316006
rect 322676 4418 322704 335326
rect 322664 4412 322716 4418
rect 322664 4354 322716 4360
rect 322112 3528 322164 3534
rect 322112 3470 322164 3476
rect 322296 3528 322348 3534
rect 322296 3470 322348 3476
rect 321468 2984 321520 2990
rect 321468 2926 321520 2932
rect 322124 480 322152 3470
rect 322768 3058 322796 336670
rect 322860 336054 322888 338014
rect 322848 336048 322900 336054
rect 322848 335990 322900 335996
rect 323228 335986 323256 338014
rect 323216 335980 323268 335986
rect 323216 335922 323268 335928
rect 322848 335504 322900 335510
rect 322848 335446 322900 335452
rect 322860 3126 322888 335446
rect 323504 325694 323532 338014
rect 323780 330478 323808 338014
rect 323872 338014 323932 338042
rect 324056 338014 324208 338042
rect 324576 338014 324728 338042
rect 324852 338014 325004 338042
rect 325128 338014 325280 338042
rect 323872 336734 323900 338014
rect 323860 336728 323912 336734
rect 323860 336670 323912 336676
rect 324056 330562 324084 338014
rect 324228 336728 324280 336734
rect 324228 336670 324280 336676
rect 324136 335980 324188 335986
rect 324136 335922 324188 335928
rect 323964 330534 324084 330562
rect 323768 330472 323820 330478
rect 323768 330414 323820 330420
rect 323504 325666 323900 325694
rect 323872 4486 323900 325666
rect 323964 4554 323992 330534
rect 324044 330472 324096 330478
rect 324044 330414 324096 330420
rect 323952 4548 324004 4554
rect 323952 4490 324004 4496
rect 323860 4480 323912 4486
rect 323860 4422 323912 4428
rect 323308 3528 323360 3534
rect 323308 3470 323360 3476
rect 322848 3120 322900 3126
rect 322848 3062 322900 3068
rect 322756 3052 322808 3058
rect 322756 2994 322808 3000
rect 323320 480 323348 3470
rect 324056 3262 324084 330414
rect 324044 3256 324096 3262
rect 324044 3198 324096 3204
rect 324148 3194 324176 335922
rect 324240 3398 324268 336670
rect 324700 336666 324728 338014
rect 324688 336660 324740 336666
rect 324688 336602 324740 336608
rect 324976 336598 325004 338014
rect 325252 336734 325280 338014
rect 325390 337770 325418 338028
rect 325772 338014 325924 338042
rect 326048 338014 326200 338042
rect 326324 338014 326476 338042
rect 325390 337742 325464 337770
rect 325240 336728 325292 336734
rect 325240 336670 325292 336676
rect 325332 336660 325384 336666
rect 325332 336602 325384 336608
rect 324964 336592 325016 336598
rect 324964 336534 325016 336540
rect 324964 336252 325016 336258
rect 324964 336194 325016 336200
rect 324976 4010 325004 336194
rect 325344 4622 325372 336602
rect 325436 4758 325464 337742
rect 325516 336728 325568 336734
rect 325516 336670 325568 336676
rect 325424 4752 325476 4758
rect 325424 4694 325476 4700
rect 325528 4690 325556 336670
rect 325896 336598 325924 338014
rect 325608 336592 325660 336598
rect 325608 336534 325660 336540
rect 325884 336592 325936 336598
rect 325884 336534 325936 336540
rect 325516 4684 325568 4690
rect 325516 4626 325568 4632
rect 325332 4616 325384 4622
rect 325332 4558 325384 4564
rect 324964 4004 325016 4010
rect 324964 3946 325016 3952
rect 325516 3596 325568 3602
rect 325516 3538 325568 3544
rect 324228 3392 324280 3398
rect 324228 3334 324280 3340
rect 324136 3188 324188 3194
rect 324136 3130 324188 3136
rect 324412 2916 324464 2922
rect 324412 2858 324464 2864
rect 324424 480 324452 2858
rect 325528 2666 325556 3538
rect 325620 2854 325648 336534
rect 326172 330478 326200 338014
rect 326448 336666 326476 338014
rect 326540 338014 326600 338042
rect 326724 338014 326968 338042
rect 327244 338014 327396 338042
rect 327520 338014 327672 338042
rect 327796 338014 328040 338042
rect 326436 336660 326488 336666
rect 326436 336602 326488 336608
rect 326540 335442 326568 338014
rect 326528 335436 326580 335442
rect 326528 335378 326580 335384
rect 326724 330562 326752 338014
rect 326804 336660 326856 336666
rect 326804 336602 326856 336608
rect 326632 330534 326752 330562
rect 326160 330472 326212 330478
rect 326160 330414 326212 330420
rect 326632 5302 326660 330534
rect 326712 330472 326764 330478
rect 326712 330414 326764 330420
rect 326724 5506 326752 330414
rect 326712 5500 326764 5506
rect 326712 5442 326764 5448
rect 326816 5438 326844 336602
rect 326988 336592 327040 336598
rect 326988 336534 327040 336540
rect 326896 335436 326948 335442
rect 326896 335378 326948 335384
rect 326804 5432 326856 5438
rect 326804 5374 326856 5380
rect 326620 5296 326672 5302
rect 326620 5238 326672 5244
rect 326804 3868 326856 3874
rect 326804 3810 326856 3816
rect 325608 2848 325660 2854
rect 325608 2790 325660 2796
rect 325528 2638 325648 2666
rect 325620 480 325648 2638
rect 326816 480 326844 3810
rect 326908 2922 326936 335378
rect 327000 3942 327028 336534
rect 327368 335850 327396 338014
rect 327644 336734 327672 338014
rect 327632 336728 327684 336734
rect 327632 336670 327684 336676
rect 327356 335844 327408 335850
rect 327356 335786 327408 335792
rect 327724 335504 327776 335510
rect 327724 335446 327776 335452
rect 326988 3936 327040 3942
rect 326988 3878 327040 3884
rect 327736 3602 327764 335446
rect 328012 5234 328040 338014
rect 328150 337770 328178 338028
rect 328380 338014 328440 338042
rect 328716 338014 328868 338042
rect 328992 338014 329236 338042
rect 329360 338014 329512 338042
rect 328150 337742 328224 337770
rect 328092 335844 328144 335850
rect 328092 335786 328144 335792
rect 328104 5370 328132 335786
rect 328092 5364 328144 5370
rect 328092 5306 328144 5312
rect 328000 5228 328052 5234
rect 328000 5170 328052 5176
rect 328196 5166 328224 337742
rect 328276 336728 328328 336734
rect 328276 336670 328328 336676
rect 328184 5160 328236 5166
rect 328184 5102 328236 5108
rect 328288 3874 328316 336670
rect 328380 4146 328408 338014
rect 328840 336666 328868 338014
rect 328828 336660 328880 336666
rect 328828 336602 328880 336608
rect 329208 335354 329236 338014
rect 329484 336734 329512 338014
rect 329576 338014 329636 338042
rect 329912 338014 330064 338042
rect 330188 338014 330432 338042
rect 330556 338014 330708 338042
rect 329472 336728 329524 336734
rect 329472 336670 329524 336676
rect 329208 335326 329512 335354
rect 329484 5030 329512 335326
rect 329472 5024 329524 5030
rect 329472 4966 329524 4972
rect 329576 4962 329604 338014
rect 329748 336728 329800 336734
rect 329748 336670 329800 336676
rect 329656 336660 329708 336666
rect 329656 336602 329708 336608
rect 329668 5098 329696 336602
rect 329656 5092 329708 5098
rect 329656 5034 329708 5040
rect 329564 4956 329616 4962
rect 329564 4898 329616 4904
rect 328368 4140 328420 4146
rect 328368 4082 328420 4088
rect 328276 3868 328328 3874
rect 328276 3810 328328 3816
rect 327724 3596 327776 3602
rect 327724 3538 327776 3544
rect 328000 3528 328052 3534
rect 328000 3470 328052 3476
rect 326896 2916 326948 2922
rect 326896 2858 326948 2864
rect 328012 480 328040 3470
rect 329196 3460 329248 3466
rect 329196 3402 329248 3408
rect 329208 480 329236 3402
rect 329760 3330 329788 336670
rect 330036 336666 330064 338014
rect 330024 336660 330076 336666
rect 330024 336602 330076 336608
rect 330404 335714 330432 338014
rect 330680 336734 330708 338014
rect 330772 338014 330832 338042
rect 331048 338014 331108 338042
rect 331384 338014 331628 338042
rect 331752 338014 331904 338042
rect 330668 336728 330720 336734
rect 330668 336670 330720 336676
rect 330392 335708 330444 335714
rect 330392 335650 330444 335656
rect 330772 4826 330800 338014
rect 330852 336728 330904 336734
rect 330852 336670 330904 336676
rect 330864 4894 330892 336670
rect 330944 336660 330996 336666
rect 330944 336602 330996 336608
rect 330852 4888 330904 4894
rect 330852 4830 330904 4836
rect 330760 4820 330812 4826
rect 330760 4762 330812 4768
rect 330392 3800 330444 3806
rect 330392 3742 330444 3748
rect 329748 3324 329800 3330
rect 329748 3266 329800 3272
rect 330404 480 330432 3742
rect 330956 3466 330984 336602
rect 331048 3534 331076 338014
rect 331600 335714 331628 338014
rect 331876 336734 331904 338014
rect 331968 338014 332028 338042
rect 332152 338014 332304 338042
rect 332428 338014 332580 338042
rect 332948 338014 333100 338042
rect 333224 338014 333376 338042
rect 333500 338014 333744 338042
rect 331864 336728 331916 336734
rect 331864 336670 331916 336676
rect 331968 336666 331996 338014
rect 331956 336660 332008 336666
rect 331956 336602 332008 336608
rect 331128 335708 331180 335714
rect 331128 335650 331180 335656
rect 331588 335708 331640 335714
rect 331588 335650 331640 335656
rect 331140 3942 331168 335650
rect 332152 9722 332180 338014
rect 332324 336728 332376 336734
rect 332324 336670 332376 336676
rect 332232 335708 332284 335714
rect 332232 335650 332284 335656
rect 332244 330585 332272 335650
rect 332230 330576 332286 330585
rect 332230 330511 332286 330520
rect 332232 330472 332284 330478
rect 332232 330414 332284 330420
rect 332140 9716 332192 9722
rect 332140 9658 332192 9664
rect 332244 7002 332272 330414
rect 332232 6996 332284 7002
rect 332232 6938 332284 6944
rect 332336 6866 332364 336670
rect 332428 330682 332456 338014
rect 332508 336660 332560 336666
rect 332508 336602 332560 336608
rect 332416 330676 332468 330682
rect 332416 330618 332468 330624
rect 332414 330576 332470 330585
rect 332414 330511 332470 330520
rect 332324 6860 332376 6866
rect 332324 6802 332376 6808
rect 332428 4214 332456 330511
rect 332416 4208 332468 4214
rect 332416 4150 332468 4156
rect 332520 4146 332548 336602
rect 333072 335850 333100 338014
rect 333060 335844 333112 335850
rect 333060 335786 333112 335792
rect 333348 335354 333376 338014
rect 333348 335326 333652 335354
rect 333624 9790 333652 335326
rect 333716 9858 333744 338014
rect 333808 338014 333868 338042
rect 334144 338014 334296 338042
rect 334420 338014 334572 338042
rect 334696 338014 334940 338042
rect 333704 9852 333756 9858
rect 333704 9794 333756 9800
rect 333612 9784 333664 9790
rect 333612 9726 333664 9732
rect 333808 6914 333836 338014
rect 334268 336666 334296 338014
rect 334256 336660 334308 336666
rect 334256 336602 334308 336608
rect 334440 336320 334492 336326
rect 334440 336262 334492 336268
rect 333888 335844 333940 335850
rect 333888 335786 333940 335792
rect 333716 6886 333836 6914
rect 332508 4140 332560 4146
rect 332508 4082 332560 4088
rect 332692 4004 332744 4010
rect 332692 3946 332744 3952
rect 331128 3936 331180 3942
rect 331128 3878 331180 3884
rect 331588 3596 331640 3602
rect 331588 3538 331640 3544
rect 331036 3528 331088 3534
rect 331036 3470 331088 3476
rect 330944 3460 330996 3466
rect 330944 3402 330996 3408
rect 331600 480 331628 3538
rect 332704 480 332732 3946
rect 333716 3738 333744 6886
rect 333900 5386 333928 335786
rect 334452 16574 334480 336262
rect 334544 325694 334572 338014
rect 334912 336734 334940 338014
rect 335004 338014 335064 338042
rect 335188 338014 335340 338042
rect 335556 338014 335616 338042
rect 335892 338014 336136 338042
rect 336260 338014 336412 338042
rect 336536 338014 336688 338042
rect 336812 338014 336964 338042
rect 337088 338014 337332 338042
rect 337456 338014 337608 338042
rect 337732 338014 337884 338042
rect 334900 336728 334952 336734
rect 334900 336670 334952 336676
rect 334544 325666 334940 325694
rect 334452 16546 334664 16574
rect 333808 5358 333928 5386
rect 333808 3874 333836 5358
rect 333888 4072 333940 4078
rect 333888 4014 333940 4020
rect 333796 3868 333848 3874
rect 333796 3810 333848 3816
rect 333704 3732 333756 3738
rect 333704 3674 333756 3680
rect 333900 480 333928 4014
rect 334636 490 334664 16546
rect 334912 9994 334940 325666
rect 335004 10062 335032 338014
rect 335084 336660 335136 336666
rect 335084 336602 335136 336608
rect 334992 10056 335044 10062
rect 334992 9998 335044 10004
rect 334900 9988 334952 9994
rect 334900 9930 334952 9936
rect 335096 9926 335124 336602
rect 335084 9920 335136 9926
rect 335084 9862 335136 9868
rect 335188 8362 335216 338014
rect 335268 336728 335320 336734
rect 335268 336670 335320 336676
rect 335176 8356 335228 8362
rect 335176 8298 335228 8304
rect 335280 4049 335308 336670
rect 335556 335782 335584 338014
rect 335728 336388 335780 336394
rect 335728 336330 335780 336336
rect 335544 335776 335596 335782
rect 335544 335718 335596 335724
rect 335740 16574 335768 336330
rect 336108 335442 336136 338014
rect 336096 335436 336148 335442
rect 336096 335378 336148 335384
rect 335740 16546 336320 16574
rect 335266 4040 335322 4049
rect 335266 3975 335322 3984
rect 334912 598 335124 626
rect 334912 490 334940 598
rect 318494 -960 318606 480
rect 319690 -960 319802 480
rect 320886 -960 320998 480
rect 322082 -960 322194 480
rect 323278 -960 323390 480
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326774 -960 326886 480
rect 327970 -960 328082 480
rect 329166 -960 329278 480
rect 330362 -960 330474 480
rect 331558 -960 331670 480
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 334636 462 334940 490
rect 335096 480 335124 598
rect 336292 480 336320 16546
rect 336384 8430 336412 338014
rect 336556 335776 336608 335782
rect 336556 335718 336608 335724
rect 336464 335436 336516 335442
rect 336464 335378 336516 335384
rect 336372 8424 336424 8430
rect 336372 8366 336424 8372
rect 336476 5574 336504 335378
rect 336464 5568 336516 5574
rect 336464 5510 336516 5516
rect 336568 3913 336596 335718
rect 336554 3904 336610 3913
rect 336554 3839 336610 3848
rect 336660 3777 336688 338014
rect 336936 335714 336964 338014
rect 337304 335986 337332 338014
rect 337580 336598 337608 338014
rect 337660 336728 337712 336734
rect 337660 336670 337712 336676
rect 337856 336682 337884 338014
rect 337948 338014 338008 338042
rect 338284 338014 338528 338042
rect 338652 338014 338804 338042
rect 338928 338014 339080 338042
rect 337948 336802 337976 338014
rect 337936 336796 337988 336802
rect 337936 336738 337988 336744
rect 337568 336592 337620 336598
rect 337568 336534 337620 336540
rect 337292 335980 337344 335986
rect 337292 335922 337344 335928
rect 336924 335708 336976 335714
rect 336924 335650 336976 335656
rect 337672 325694 337700 336670
rect 337856 336654 338068 336682
rect 337752 335980 337804 335986
rect 337752 335922 337804 335928
rect 337764 330562 337792 335922
rect 337936 335708 337988 335714
rect 337936 335650 337988 335656
rect 337764 330534 337884 330562
rect 337672 325666 337792 325694
rect 337764 8566 337792 325666
rect 337752 8560 337804 8566
rect 337752 8502 337804 8508
rect 337856 8498 337884 330534
rect 337844 8492 337896 8498
rect 337844 8434 337896 8440
rect 337948 5642 337976 335650
rect 338040 5710 338068 336654
rect 338500 335850 338528 338014
rect 338776 336734 338804 338014
rect 338764 336728 338816 336734
rect 338764 336670 338816 336676
rect 338764 336592 338816 336598
rect 338764 336534 338816 336540
rect 338580 336184 338632 336190
rect 338580 336126 338632 336132
rect 338488 335844 338540 335850
rect 338488 335786 338540 335792
rect 338592 16574 338620 336126
rect 338592 16546 338712 16574
rect 338028 5704 338080 5710
rect 338028 5646 338080 5652
rect 337936 5636 337988 5642
rect 337936 5578 337988 5584
rect 336646 3768 336702 3777
rect 336646 3703 336702 3712
rect 337476 3664 337528 3670
rect 337476 3606 337528 3612
rect 337488 480 337516 3606
rect 338684 480 338712 16546
rect 338776 3670 338804 336534
rect 339052 325694 339080 338014
rect 339190 337770 339218 338028
rect 339328 338014 339480 338042
rect 339848 338014 340000 338042
rect 340124 338014 340276 338042
rect 340400 338014 340552 338042
rect 339190 337742 339264 337770
rect 339236 336734 339264 337742
rect 339132 336728 339184 336734
rect 339132 336670 339184 336676
rect 339224 336728 339276 336734
rect 339224 336670 339276 336676
rect 339144 330562 339172 336670
rect 339144 330534 339264 330562
rect 339052 325666 339172 325694
rect 339144 8634 339172 325666
rect 339132 8628 339184 8634
rect 339132 8570 339184 8576
rect 339236 5778 339264 330534
rect 339328 5846 339356 338014
rect 339408 336728 339460 336734
rect 339408 336670 339460 336676
rect 339316 5840 339368 5846
rect 339316 5782 339368 5788
rect 339224 5772 339276 5778
rect 339224 5714 339276 5720
rect 338764 3664 338816 3670
rect 339420 3641 339448 336670
rect 339972 336666 340000 338014
rect 339960 336660 340012 336666
rect 339960 336602 340012 336608
rect 339868 336116 339920 336122
rect 339868 336058 339920 336064
rect 338764 3606 338816 3612
rect 339406 3632 339462 3641
rect 339406 3567 339462 3576
rect 339880 480 339908 336058
rect 340248 335918 340276 338014
rect 340524 336734 340552 338014
rect 340616 338014 340676 338042
rect 341044 338014 341196 338042
rect 341320 338014 341472 338042
rect 341596 338014 341748 338042
rect 341872 338014 342024 338042
rect 340512 336728 340564 336734
rect 340512 336670 340564 336676
rect 340236 335912 340288 335918
rect 340236 335854 340288 335860
rect 340616 8770 340644 338014
rect 340788 336728 340840 336734
rect 340788 336670 340840 336676
rect 340696 336660 340748 336666
rect 340696 336602 340748 336608
rect 340604 8764 340656 8770
rect 340604 8706 340656 8712
rect 340708 8702 340736 336602
rect 340696 8696 340748 8702
rect 340696 8638 340748 8644
rect 340800 5914 340828 336670
rect 341168 336598 341196 338014
rect 341444 336734 341472 338014
rect 341432 336728 341484 336734
rect 341432 336670 341484 336676
rect 341156 336592 341208 336598
rect 341156 336534 341208 336540
rect 341720 335354 341748 338014
rect 341996 336530 342024 338014
rect 342088 338014 342240 338042
rect 342516 338014 342668 338042
rect 342792 338014 342944 338042
rect 343068 338014 343220 338042
rect 341984 336524 342036 336530
rect 341984 336466 342036 336472
rect 341720 335326 342024 335354
rect 341996 8838 342024 335326
rect 341984 8832 342036 8838
rect 341984 8774 342036 8780
rect 342088 6050 342116 338014
rect 342640 336734 342668 338014
rect 342168 336728 342220 336734
rect 342168 336670 342220 336676
rect 342628 336728 342680 336734
rect 342628 336670 342680 336676
rect 342076 6044 342128 6050
rect 342076 5986 342128 5992
rect 342180 5982 342208 336670
rect 342916 336666 342944 338014
rect 342904 336660 342956 336666
rect 342904 336602 342956 336608
rect 343192 335986 343220 338014
rect 343284 338014 343436 338042
rect 343712 338014 343864 338042
rect 343988 338014 344140 338042
rect 344264 338014 344508 338042
rect 344632 338014 344784 338042
rect 343180 335980 343232 335986
rect 343180 335922 343232 335928
rect 343284 9654 343312 338014
rect 343364 336728 343416 336734
rect 343364 336670 343416 336676
rect 343272 9648 343324 9654
rect 343272 9590 343324 9596
rect 343376 8906 343404 336670
rect 343836 336666 343864 338014
rect 343548 336660 343600 336666
rect 343548 336602 343600 336608
rect 343824 336660 343876 336666
rect 343824 336602 343876 336608
rect 343456 335980 343508 335986
rect 343456 335922 343508 335928
rect 343364 8900 343416 8906
rect 343364 8842 343416 8848
rect 343468 6118 343496 335922
rect 343456 6112 343508 6118
rect 343456 6054 343508 6060
rect 342168 5976 342220 5982
rect 342168 5918 342220 5924
rect 340788 5908 340840 5914
rect 340788 5850 340840 5856
rect 343560 3806 343588 336602
rect 344112 336326 344140 338014
rect 344100 336320 344152 336326
rect 344100 336262 344152 336268
rect 344480 335354 344508 338014
rect 344756 336462 344784 338014
rect 344848 338014 344908 338042
rect 345184 338014 345336 338042
rect 345460 338014 345704 338042
rect 345828 338014 345980 338042
rect 344744 336456 344796 336462
rect 344744 336398 344796 336404
rect 344744 336320 344796 336326
rect 344744 336262 344796 336268
rect 344480 335326 344692 335354
rect 344664 9586 344692 335326
rect 344652 9580 344704 9586
rect 344652 9522 344704 9528
rect 344756 6798 344784 336262
rect 344744 6792 344796 6798
rect 344744 6734 344796 6740
rect 344848 6730 344876 338014
rect 345308 336666 345336 338014
rect 344928 336660 344980 336666
rect 344928 336602 344980 336608
rect 345296 336660 345348 336666
rect 345296 336602 345348 336608
rect 344836 6724 344888 6730
rect 344836 6666 344888 6672
rect 342168 3800 342220 3806
rect 342168 3742 342220 3748
rect 343548 3800 343600 3806
rect 343548 3742 343600 3748
rect 340972 2984 341024 2990
rect 340972 2926 341024 2932
rect 340984 480 341012 2926
rect 342180 480 342208 3742
rect 344560 3120 344612 3126
rect 344560 3062 344612 3068
rect 343364 3052 343416 3058
rect 343364 2994 343416 3000
rect 343376 480 343404 2994
rect 344572 480 344600 3062
rect 344940 2990 344968 336602
rect 345676 336394 345704 338014
rect 345952 336598 345980 338014
rect 346090 337770 346118 338028
rect 346320 338014 346380 338042
rect 346656 338014 346900 338042
rect 347024 338014 347176 338042
rect 347300 338014 347452 338042
rect 346090 337742 346164 337770
rect 346032 336660 346084 336666
rect 346032 336602 346084 336608
rect 345940 336592 345992 336598
rect 345940 336534 345992 336540
rect 345664 336388 345716 336394
rect 345664 336330 345716 336336
rect 346044 9518 346072 336602
rect 346032 9512 346084 9518
rect 346032 9454 346084 9460
rect 346136 9450 346164 337742
rect 346216 336592 346268 336598
rect 346216 336534 346268 336540
rect 346320 336546 346348 338014
rect 346872 336666 346900 338014
rect 346860 336660 346912 336666
rect 346860 336602 346912 336608
rect 346124 9444 346176 9450
rect 346124 9386 346176 9392
rect 346228 6662 346256 336534
rect 346320 336518 346440 336546
rect 346308 336388 346360 336394
rect 346308 336330 346360 336336
rect 346216 6656 346268 6662
rect 346216 6598 346268 6604
rect 345756 4412 345808 4418
rect 345756 4354 345808 4360
rect 344928 2984 344980 2990
rect 344928 2926 344980 2932
rect 345768 480 345796 4354
rect 346320 3058 346348 336330
rect 346412 336190 346440 336518
rect 346400 336184 346452 336190
rect 346400 336126 346452 336132
rect 346768 336048 346820 336054
rect 346768 335990 346820 335996
rect 346780 16574 346808 335990
rect 347148 325694 347176 338014
rect 347424 336598 347452 338014
rect 347562 337770 347590 338028
rect 347852 338014 348096 338042
rect 348220 338014 348372 338042
rect 348496 338014 348648 338042
rect 348772 338014 348924 338042
rect 347562 337742 347636 337770
rect 347504 336660 347556 336666
rect 347504 336602 347556 336608
rect 347412 336592 347464 336598
rect 347412 336534 347464 336540
rect 347148 325666 347452 325694
rect 346780 16546 346992 16574
rect 346308 3052 346360 3058
rect 346308 2994 346360 3000
rect 346964 480 346992 16546
rect 347424 9382 347452 325666
rect 347412 9376 347464 9382
rect 347412 9318 347464 9324
rect 347516 6594 347544 336602
rect 347504 6588 347556 6594
rect 347504 6530 347556 6536
rect 347608 6526 347636 337742
rect 348068 336598 348096 338014
rect 347688 336592 347740 336598
rect 347688 336534 347740 336540
rect 348056 336592 348108 336598
rect 348056 336534 348108 336540
rect 347596 6520 347648 6526
rect 347596 6462 347648 6468
rect 347700 3126 347728 336534
rect 348344 336122 348372 338014
rect 348620 336666 348648 338014
rect 348896 336682 348924 338014
rect 349034 337770 349062 338028
rect 349416 338014 349568 338042
rect 349692 338014 349844 338042
rect 349968 338014 350120 338042
rect 350244 338014 350396 338042
rect 350612 338014 350764 338042
rect 350888 338014 351040 338042
rect 351164 338014 351316 338042
rect 351440 338014 351684 338042
rect 349034 337742 349108 337770
rect 349080 336818 349108 337742
rect 349080 336790 349200 336818
rect 348608 336660 348660 336666
rect 348896 336654 349016 336682
rect 348608 336602 348660 336608
rect 348884 336592 348936 336598
rect 348884 336534 348936 336540
rect 348332 336116 348384 336122
rect 348332 336058 348384 336064
rect 348896 9314 348924 336534
rect 348884 9308 348936 9314
rect 348884 9250 348936 9256
rect 348988 9246 349016 336654
rect 349068 336660 349120 336666
rect 349068 336602 349120 336608
rect 348976 9240 349028 9246
rect 348976 9182 349028 9188
rect 349080 6458 349108 336602
rect 349172 336326 349200 336790
rect 349540 336598 349568 338014
rect 349816 336666 349844 338014
rect 349804 336660 349856 336666
rect 349804 336602 349856 336608
rect 349528 336592 349580 336598
rect 349528 336534 349580 336540
rect 349160 336320 349212 336326
rect 349160 336262 349212 336268
rect 350092 336258 350120 338014
rect 350264 336660 350316 336666
rect 350264 336602 350316 336608
rect 350080 336252 350132 336258
rect 350080 336194 350132 336200
rect 350276 9178 350304 336602
rect 350264 9172 350316 9178
rect 350264 9114 350316 9120
rect 349068 6452 349120 6458
rect 349068 6394 349120 6400
rect 350368 6322 350396 338014
rect 350736 336598 350764 338014
rect 350448 336592 350500 336598
rect 350448 336534 350500 336540
rect 350724 336592 350776 336598
rect 350724 336534 350776 336540
rect 350460 6390 350488 336534
rect 351012 336394 351040 338014
rect 351288 336666 351316 338014
rect 351276 336660 351328 336666
rect 351276 336602 351328 336608
rect 351552 336592 351604 336598
rect 351552 336534 351604 336540
rect 351000 336388 351052 336394
rect 351000 336330 351052 336336
rect 351564 9110 351592 336534
rect 351552 9104 351604 9110
rect 351552 9046 351604 9052
rect 351656 9042 351684 338014
rect 351794 337770 351822 338028
rect 352084 338014 352236 338042
rect 352360 338014 352512 338042
rect 352636 338014 352880 338042
rect 351794 337742 351868 337770
rect 351736 336660 351788 336666
rect 351736 336602 351788 336608
rect 351644 9036 351696 9042
rect 351644 8978 351696 8984
rect 350448 6384 350500 6390
rect 350448 6326 350500 6332
rect 350356 6316 350408 6322
rect 350356 6258 350408 6264
rect 351748 6254 351776 336602
rect 351840 336546 351868 337742
rect 351840 336518 351960 336546
rect 351828 336388 351880 336394
rect 351828 336330 351880 336336
rect 351736 6248 351788 6254
rect 351736 6190 351788 6196
rect 349252 4480 349304 4486
rect 349252 4422 349304 4428
rect 348056 3188 348108 3194
rect 348056 3130 348108 3136
rect 347688 3120 347740 3126
rect 347688 3062 347740 3068
rect 348068 480 348096 3130
rect 349264 480 349292 4422
rect 351644 3392 351696 3398
rect 351644 3334 351696 3340
rect 350448 3256 350500 3262
rect 350448 3198 350500 3204
rect 350460 480 350488 3198
rect 351656 480 351684 3334
rect 351840 3194 351868 336330
rect 351932 336190 351960 336518
rect 351920 336184 351972 336190
rect 351920 336126 351972 336132
rect 352208 335374 352236 338014
rect 352196 335368 352248 335374
rect 352196 335310 352248 335316
rect 352484 325694 352512 338014
rect 352852 336326 352880 338014
rect 352990 337770 353018 338028
rect 353128 338014 353280 338042
rect 353556 338014 353708 338042
rect 353832 338014 354076 338042
rect 354200 338014 354352 338042
rect 354476 338014 354628 338042
rect 354752 338014 354904 338042
rect 355028 338014 355272 338042
rect 355396 338014 355548 338042
rect 355672 338014 355824 338042
rect 352990 337742 353064 337770
rect 352932 336660 352984 336666
rect 352932 336602 352984 336608
rect 352840 336320 352892 336326
rect 352840 336262 352892 336268
rect 352484 325666 352880 325694
rect 352852 8974 352880 325666
rect 352944 9217 352972 336602
rect 352930 9208 352986 9217
rect 352930 9143 352986 9152
rect 352840 8968 352892 8974
rect 352840 8910 352892 8916
rect 353036 6633 353064 337742
rect 353128 336666 353156 338014
rect 353116 336660 353168 336666
rect 353116 336602 353168 336608
rect 353208 336320 353260 336326
rect 353208 336262 353260 336268
rect 353116 335232 353168 335238
rect 353116 335174 353168 335180
rect 353022 6624 353078 6633
rect 353022 6559 353078 6568
rect 353128 6186 353156 335174
rect 353116 6180 353168 6186
rect 353116 6122 353168 6128
rect 352840 4548 352892 4554
rect 352840 4490 352892 4496
rect 351828 3188 351880 3194
rect 351828 3130 351880 3136
rect 352852 480 352880 4490
rect 353220 3262 353248 336262
rect 353680 336122 353708 338014
rect 354048 336666 354076 338014
rect 354036 336660 354088 336666
rect 354036 336602 354088 336608
rect 353668 336116 353720 336122
rect 353668 336058 353720 336064
rect 354324 335354 354352 338014
rect 354496 336660 354548 336666
rect 354496 336602 354548 336608
rect 354324 335326 354444 335354
rect 354416 9081 354444 335326
rect 354402 9072 354458 9081
rect 354402 9007 354458 9016
rect 354508 6497 354536 336602
rect 354494 6488 354550 6497
rect 354494 6423 354550 6432
rect 354036 4616 354088 4622
rect 354036 4558 354088 4564
rect 353208 3256 353260 3262
rect 353208 3198 353260 3204
rect 354048 480 354076 4558
rect 354600 3398 354628 338014
rect 354876 336598 354904 338014
rect 354864 336592 354916 336598
rect 354864 336534 354916 336540
rect 355244 335714 355272 338014
rect 355232 335708 355284 335714
rect 355232 335650 355284 335656
rect 355520 335646 355548 338014
rect 355692 336592 355744 336598
rect 355692 336534 355744 336540
rect 355508 335640 355560 335646
rect 355508 335582 355560 335588
rect 355704 10198 355732 336534
rect 355796 10266 355824 338014
rect 355934 337770 355962 338028
rect 356224 338014 356468 338042
rect 356592 338014 356744 338042
rect 356868 338014 357020 338042
rect 357144 338014 357296 338042
rect 355934 337742 356008 337770
rect 355876 335708 355928 335714
rect 355876 335650 355928 335656
rect 355784 10260 355836 10266
rect 355784 10202 355836 10208
rect 355692 10192 355744 10198
rect 355692 10134 355744 10140
rect 355888 10130 355916 335650
rect 355876 10124 355928 10130
rect 355876 10066 355928 10072
rect 355980 8945 356008 337742
rect 356440 335782 356468 338014
rect 356428 335776 356480 335782
rect 356428 335718 356480 335724
rect 356716 335354 356744 338014
rect 356992 336682 357020 338014
rect 356992 336654 357204 336682
rect 356716 335326 357112 335354
rect 357084 11014 357112 335326
rect 357176 330562 357204 336654
rect 357268 330698 357296 338014
rect 357360 338014 357420 338042
rect 357788 338014 357940 338042
rect 358064 338014 358216 338042
rect 358340 338014 358492 338042
rect 357360 330834 357388 338014
rect 357912 336054 357940 338014
rect 357900 336048 357952 336054
rect 357900 335990 357952 335996
rect 358188 335354 358216 338014
rect 358464 336682 358492 338014
rect 358602 337770 358630 338028
rect 358984 338014 359136 338042
rect 359260 338014 359412 338042
rect 359536 338014 359688 338042
rect 358602 337742 358676 337770
rect 358464 336654 358584 336682
rect 358188 335326 358492 335354
rect 357360 330806 357480 330834
rect 357268 330670 357388 330698
rect 357176 330534 357296 330562
rect 357164 330472 357216 330478
rect 357164 330414 357216 330420
rect 357072 11008 357124 11014
rect 357072 10950 357124 10956
rect 357176 10742 357204 330414
rect 357268 10878 357296 330534
rect 357360 10946 357388 330670
rect 357452 330478 357480 330806
rect 357440 330472 357492 330478
rect 357440 330414 357492 330420
rect 357348 10940 357400 10946
rect 357348 10882 357400 10888
rect 357256 10872 357308 10878
rect 357256 10814 357308 10820
rect 357164 10736 357216 10742
rect 357164 10678 357216 10684
rect 358464 10674 358492 335326
rect 358452 10668 358504 10674
rect 358452 10610 358504 10616
rect 358556 10606 358584 336654
rect 358544 10600 358596 10606
rect 358544 10542 358596 10548
rect 358648 10538 358676 337742
rect 359108 336054 359136 338014
rect 358728 336048 358780 336054
rect 358728 335990 358780 335996
rect 359096 336048 359148 336054
rect 359096 335990 359148 335996
rect 358740 10810 358768 335990
rect 359384 325694 359412 338014
rect 359660 336598 359688 338014
rect 359798 337770 359826 338028
rect 360028 338014 360180 338042
rect 360456 338014 360608 338042
rect 360732 338014 360884 338042
rect 361008 338014 361252 338042
rect 359798 337742 359872 337770
rect 359648 336592 359700 336598
rect 359648 336534 359700 336540
rect 359384 325666 359780 325694
rect 358728 10804 358780 10810
rect 358728 10746 358780 10752
rect 358636 10532 358688 10538
rect 358636 10474 358688 10480
rect 359752 10402 359780 325666
rect 359740 10396 359792 10402
rect 359740 10338 359792 10344
rect 359844 10334 359872 337742
rect 359924 336048 359976 336054
rect 359924 335990 359976 335996
rect 359936 10470 359964 335990
rect 360028 10577 360056 338014
rect 360580 336598 360608 338014
rect 360108 336592 360160 336598
rect 360108 336534 360160 336540
rect 360568 336592 360620 336598
rect 360568 336534 360620 336540
rect 360014 10568 360070 10577
rect 360014 10503 360070 10512
rect 359924 10464 359976 10470
rect 359924 10406 359976 10412
rect 359832 10328 359884 10334
rect 359832 10270 359884 10276
rect 355966 8936 356022 8945
rect 355966 8871 356022 8880
rect 360120 7070 360148 336534
rect 360856 325694 360884 338014
rect 361224 335714 361252 338014
rect 361362 337770 361390 338028
rect 361652 338014 361804 338042
rect 361928 338014 362080 338042
rect 362204 338014 362448 338042
rect 361362 337742 361436 337770
rect 361304 336592 361356 336598
rect 361304 336534 361356 336540
rect 361212 335708 361264 335714
rect 361212 335650 361264 335656
rect 360856 325666 361252 325694
rect 361224 10441 361252 325666
rect 361210 10432 361266 10441
rect 361210 10367 361266 10376
rect 361316 7138 361344 336534
rect 361408 7206 361436 337742
rect 361776 336054 361804 338014
rect 361764 336048 361816 336054
rect 361764 335990 361816 335996
rect 362052 335850 362080 338014
rect 362420 336598 362448 338014
rect 362512 338014 362572 338042
rect 362788 338014 362848 338042
rect 363124 338014 363276 338042
rect 363400 338014 363644 338042
rect 363768 338014 363920 338042
rect 362408 336592 362460 336598
rect 362408 336534 362460 336540
rect 362040 335844 362092 335850
rect 362040 335786 362092 335792
rect 361488 335708 361540 335714
rect 361488 335650 361540 335656
rect 361396 7200 361448 7206
rect 361396 7142 361448 7148
rect 361304 7132 361356 7138
rect 361304 7074 361356 7080
rect 360108 7064 360160 7070
rect 360108 7006 360160 7012
rect 359924 5500 359976 5506
rect 359924 5442 359976 5448
rect 357532 4752 357584 4758
rect 357532 4694 357584 4700
rect 356336 4684 356388 4690
rect 356336 4626 356388 4632
rect 354588 3392 354640 3398
rect 354588 3334 354640 3340
rect 355232 2848 355284 2854
rect 355232 2790 355284 2796
rect 355244 480 355272 2790
rect 356348 480 356376 4626
rect 357544 480 357572 4694
rect 358728 2916 358780 2922
rect 358728 2858 358780 2864
rect 358740 480 358768 2858
rect 359936 480 359964 5442
rect 361120 5432 361172 5438
rect 361120 5374 361172 5380
rect 361132 480 361160 5374
rect 361500 4282 361528 335650
rect 362512 12238 362540 338014
rect 362684 336592 362736 336598
rect 362684 336534 362736 336540
rect 362592 336048 362644 336054
rect 362592 335990 362644 335996
rect 362500 12232 362552 12238
rect 362500 12174 362552 12180
rect 362604 10305 362632 335990
rect 362590 10296 362646 10305
rect 362590 10231 362646 10240
rect 362696 7274 362724 336534
rect 362684 7268 362736 7274
rect 362684 7210 362736 7216
rect 362788 4418 362816 338014
rect 363248 336598 363276 338014
rect 363236 336592 363288 336598
rect 363236 336534 363288 336540
rect 362868 335844 362920 335850
rect 362868 335786 362920 335792
rect 362776 4412 362828 4418
rect 362776 4354 362828 4360
rect 362880 4350 362908 335786
rect 363616 325694 363644 338014
rect 363892 335510 363920 338014
rect 364030 337770 364058 338028
rect 364260 338014 364320 338042
rect 364596 338014 364840 338042
rect 364964 338014 365116 338042
rect 365240 338014 365392 338042
rect 365516 338014 365668 338042
rect 365792 338014 366036 338042
rect 366160 338014 366312 338042
rect 366436 338014 366588 338042
rect 366712 338014 366864 338042
rect 364030 337742 364104 337770
rect 363880 335504 363932 335510
rect 363880 335446 363932 335452
rect 363616 325666 364012 325694
rect 363984 12170 364012 325666
rect 363972 12164 364024 12170
rect 363972 12106 364024 12112
rect 364076 7410 364104 337742
rect 364156 336592 364208 336598
rect 364156 336534 364208 336540
rect 364064 7404 364116 7410
rect 364064 7346 364116 7352
rect 364168 7342 364196 336534
rect 364260 335850 364288 338014
rect 364248 335844 364300 335850
rect 364248 335786 364300 335792
rect 364812 335646 364840 338014
rect 364800 335640 364852 335646
rect 364800 335582 364852 335588
rect 364248 335504 364300 335510
rect 364248 335446 364300 335452
rect 364156 7336 364208 7342
rect 364156 7278 364208 7284
rect 363512 5296 363564 5302
rect 363512 5238 363564 5244
rect 362868 4344 362920 4350
rect 362868 4286 362920 4292
rect 361488 4276 361540 4282
rect 361488 4218 361540 4224
rect 362316 3324 362368 3330
rect 362316 3266 362368 3272
rect 362328 480 362356 3266
rect 363524 480 363552 5238
rect 364260 4486 364288 335446
rect 365088 335354 365116 338014
rect 365364 335578 365392 338014
rect 365536 335640 365588 335646
rect 365536 335582 365588 335588
rect 365352 335572 365404 335578
rect 365352 335514 365404 335520
rect 365088 335326 365484 335354
rect 365456 7478 365484 335326
rect 365444 7472 365496 7478
rect 365444 7414 365496 7420
rect 364616 5364 364668 5370
rect 364616 5306 364668 5312
rect 364248 4480 364300 4486
rect 364248 4422 364300 4428
rect 364628 480 364656 5306
rect 365548 4554 365576 335582
rect 365640 4622 365668 338014
rect 366008 335714 366036 338014
rect 366284 335850 366312 338014
rect 366272 335844 366324 335850
rect 366272 335786 366324 335792
rect 366560 335782 366588 338014
rect 366732 335844 366784 335850
rect 366732 335786 366784 335792
rect 366548 335776 366600 335782
rect 366548 335718 366600 335724
rect 365996 335708 366048 335714
rect 365996 335650 366048 335656
rect 366744 12102 366772 335786
rect 366732 12096 366784 12102
rect 366732 12038 366784 12044
rect 366836 8294 366864 338014
rect 366928 338014 366988 338042
rect 367356 338014 367508 338042
rect 367632 338014 367784 338042
rect 367908 338014 368060 338042
rect 368184 338014 368428 338042
rect 368552 338014 368704 338042
rect 368828 338014 368980 338042
rect 369104 338014 369256 338042
rect 369380 338014 369624 338042
rect 366928 335850 366956 338014
rect 366916 335844 366968 335850
rect 366916 335786 366968 335792
rect 367480 335782 367508 338014
rect 367756 335850 367784 338014
rect 367744 335844 367796 335850
rect 367744 335786 367796 335792
rect 367008 335776 367060 335782
rect 367008 335718 367060 335724
rect 367468 335776 367520 335782
rect 367468 335718 367520 335724
rect 366916 335708 366968 335714
rect 366916 335650 366968 335656
rect 366824 8288 366876 8294
rect 366824 8230 366876 8236
rect 366928 7546 366956 335650
rect 366916 7540 366968 7546
rect 366916 7482 366968 7488
rect 367020 6914 367048 335718
rect 368032 335354 368060 338014
rect 368204 335844 368256 335850
rect 368204 335786 368256 335792
rect 368032 335326 368152 335354
rect 368124 12034 368152 335326
rect 368112 12028 368164 12034
rect 368112 11970 368164 11976
rect 368216 8226 368244 335786
rect 368296 335776 368348 335782
rect 368296 335718 368348 335724
rect 368204 8220 368256 8226
rect 368204 8162 368256 8168
rect 366928 6886 367048 6914
rect 366928 4690 366956 6886
rect 367008 5228 367060 5234
rect 367008 5170 367060 5176
rect 366916 4684 366968 4690
rect 366916 4626 366968 4632
rect 365628 4616 365680 4622
rect 365628 4558 365680 4564
rect 365536 4548 365588 4554
rect 365536 4490 365588 4496
rect 365812 4140 365864 4146
rect 365812 4082 365864 4088
rect 365824 480 365852 4082
rect 367020 480 367048 5170
rect 368204 5160 368256 5166
rect 368204 5102 368256 5108
rect 368216 480 368244 5102
rect 368308 4758 368336 335718
rect 368400 5506 368428 338014
rect 368676 335782 368704 338014
rect 368664 335776 368716 335782
rect 368664 335718 368716 335724
rect 368952 335646 368980 338014
rect 369228 335850 369256 338014
rect 369216 335844 369268 335850
rect 369216 335786 369268 335792
rect 369492 335776 369544 335782
rect 369492 335718 369544 335724
rect 368940 335640 368992 335646
rect 368940 335582 368992 335588
rect 369504 8158 369532 335718
rect 369492 8152 369544 8158
rect 369492 8094 369544 8100
rect 369596 8090 369624 338014
rect 369734 337770 369762 338028
rect 370024 338014 370176 338042
rect 370300 338014 370452 338042
rect 370576 338014 370820 338042
rect 370944 338014 371096 338042
rect 369734 337742 369808 337770
rect 369676 335844 369728 335850
rect 369676 335786 369728 335792
rect 369584 8084 369636 8090
rect 369584 8026 369636 8032
rect 368388 5500 368440 5506
rect 368388 5442 368440 5448
rect 369688 5438 369716 335786
rect 369676 5432 369728 5438
rect 369676 5374 369728 5380
rect 368296 4752 368348 4758
rect 368296 4694 368348 4700
rect 369780 3602 369808 337742
rect 370148 330546 370176 338014
rect 370424 335374 370452 338014
rect 370792 335850 370820 338014
rect 370780 335844 370832 335850
rect 370780 335786 370832 335792
rect 370412 335368 370464 335374
rect 370412 335310 370464 335316
rect 370872 335368 370924 335374
rect 370872 335310 370924 335316
rect 370964 335368 371016 335374
rect 370964 335310 371016 335316
rect 370136 330540 370188 330546
rect 370136 330482 370188 330488
rect 370884 8022 370912 335310
rect 370872 8016 370924 8022
rect 370872 7958 370924 7964
rect 370976 7954 371004 335310
rect 371068 331214 371096 338014
rect 371160 338014 371220 338042
rect 371496 338014 371648 338042
rect 371772 338014 372016 338042
rect 372140 338014 372292 338042
rect 372416 338014 372568 338042
rect 372692 338014 372844 338042
rect 372968 338014 373212 338042
rect 373336 338014 373488 338042
rect 371160 335374 371188 338014
rect 371620 335374 371648 338014
rect 371988 335442 372016 338014
rect 371976 335436 372028 335442
rect 371976 335378 372028 335384
rect 371148 335368 371200 335374
rect 371148 335310 371200 335316
rect 371608 335368 371660 335374
rect 371608 335310 371660 335316
rect 372160 335368 372212 335374
rect 372160 335310 372212 335316
rect 372172 331214 372200 335310
rect 372264 334642 372292 338014
rect 372540 335782 372568 338014
rect 372528 335776 372580 335782
rect 372528 335718 372580 335724
rect 372816 335442 372844 338014
rect 372528 335436 372580 335442
rect 372528 335378 372580 335384
rect 372804 335436 372856 335442
rect 372804 335378 372856 335384
rect 372264 334614 372476 334642
rect 371068 331186 371188 331214
rect 372172 331186 372384 331214
rect 371056 330540 371108 330546
rect 371056 330482 371108 330488
rect 370964 7948 371016 7954
rect 370964 7890 371016 7896
rect 371068 5370 371096 330482
rect 371056 5364 371108 5370
rect 371056 5306 371108 5312
rect 371160 5302 371188 331186
rect 372356 11966 372384 331186
rect 372344 11960 372396 11966
rect 372344 11902 372396 11908
rect 372448 7886 372476 334614
rect 372436 7880 372488 7886
rect 372436 7822 372488 7828
rect 371148 5296 371200 5302
rect 371148 5238 371200 5244
rect 372540 5234 372568 335378
rect 373184 335374 373212 338014
rect 373172 335368 373224 335374
rect 373172 335310 373224 335316
rect 373460 325694 373488 338014
rect 373598 337770 373626 338028
rect 373736 338014 373888 338042
rect 374164 338014 374408 338042
rect 374532 338014 374684 338042
rect 374808 338014 374960 338042
rect 373598 337742 373672 337770
rect 373644 335374 373672 337742
rect 373540 335368 373592 335374
rect 373540 335310 373592 335316
rect 373632 335368 373684 335374
rect 373632 335310 373684 335316
rect 373552 331214 373580 335310
rect 373552 331186 373672 331214
rect 373460 325666 373580 325694
rect 373552 11898 373580 325666
rect 373540 11892 373592 11898
rect 373540 11834 373592 11840
rect 373644 7818 373672 331186
rect 373632 7812 373684 7818
rect 373632 7754 373684 7760
rect 373736 7750 373764 338014
rect 373908 335436 373960 335442
rect 373908 335378 373960 335384
rect 373816 335368 373868 335374
rect 373816 335310 373868 335316
rect 373724 7744 373776 7750
rect 373724 7686 373776 7692
rect 372528 5228 372580 5234
rect 372528 5170 372580 5176
rect 373828 5098 373856 335310
rect 373920 5166 373948 335378
rect 374380 330546 374408 338014
rect 374656 335374 374684 338014
rect 374644 335368 374696 335374
rect 374644 335310 374696 335316
rect 374368 330540 374420 330546
rect 374368 330482 374420 330488
rect 374932 7682 374960 338014
rect 375070 337770 375098 338028
rect 375208 338014 375360 338042
rect 375728 338014 375880 338042
rect 376004 338014 376156 338042
rect 376280 338014 376432 338042
rect 375070 337742 375144 337770
rect 375116 335374 375144 337742
rect 375012 335368 375064 335374
rect 375012 335310 375064 335316
rect 375104 335368 375156 335374
rect 375104 335310 375156 335316
rect 374920 7676 374972 7682
rect 374920 7618 374972 7624
rect 373908 5160 373960 5166
rect 373908 5102 373960 5108
rect 370596 5092 370648 5098
rect 370596 5034 370648 5040
rect 373816 5092 373868 5098
rect 373816 5034 373868 5040
rect 369400 3596 369452 3602
rect 369400 3538 369452 3544
rect 369768 3596 369820 3602
rect 369768 3538 369820 3544
rect 369412 480 369440 3538
rect 370608 480 370636 5034
rect 375024 5030 375052 335310
rect 375208 331214 375236 338014
rect 375852 335374 375880 338014
rect 376128 336802 376156 338014
rect 376116 336796 376168 336802
rect 376116 336738 376168 336744
rect 375288 335368 375340 335374
rect 375288 335310 375340 335316
rect 375840 335368 375892 335374
rect 375840 335310 375892 335316
rect 375116 331186 375236 331214
rect 371700 5024 371752 5030
rect 371700 4966 371752 4972
rect 375012 5024 375064 5030
rect 375012 4966 375064 4972
rect 371712 480 371740 4966
rect 375116 4962 375144 331186
rect 375196 330540 375248 330546
rect 375196 330482 375248 330488
rect 374092 4956 374144 4962
rect 374092 4898 374144 4904
rect 375104 4956 375156 4962
rect 375104 4898 375156 4904
rect 372896 3528 372948 3534
rect 372896 3470 372948 3476
rect 372908 480 372936 3470
rect 374104 480 374132 4898
rect 375208 3534 375236 330482
rect 375300 3618 375328 335310
rect 376404 330546 376432 338014
rect 376542 337770 376570 338028
rect 376924 338014 377076 338042
rect 377200 338014 377352 338042
rect 377476 338014 377628 338042
rect 377752 338014 377904 338042
rect 376542 337742 376616 337770
rect 376484 335368 376536 335374
rect 376484 335310 376536 335316
rect 376392 330540 376444 330546
rect 376392 330482 376444 330488
rect 376496 7614 376524 335310
rect 376588 7993 376616 337742
rect 377048 335442 377076 338014
rect 377036 335436 377088 335442
rect 377036 335378 377088 335384
rect 377324 335374 377352 338014
rect 377404 335572 377456 335578
rect 377404 335514 377456 335520
rect 377312 335368 377364 335374
rect 377312 335310 377364 335316
rect 376668 330540 376720 330546
rect 376668 330482 376720 330488
rect 376574 7984 376630 7993
rect 376574 7919 376630 7928
rect 376484 7608 376536 7614
rect 376484 7550 376536 7556
rect 376680 5273 376708 330482
rect 377416 10713 377444 335514
rect 377600 331214 377628 338014
rect 377876 336433 377904 338014
rect 377968 338014 378120 338042
rect 378396 338014 378548 338042
rect 378672 338014 378824 338042
rect 378948 338014 379100 338042
rect 377862 336424 377918 336433
rect 377862 336359 377918 336368
rect 377600 331186 377904 331214
rect 377402 10704 377458 10713
rect 377402 10639 377458 10648
rect 377876 7857 377904 331186
rect 377862 7848 377918 7857
rect 377862 7783 377918 7792
rect 376666 5264 376722 5273
rect 376666 5199 376722 5208
rect 377968 5137 377996 338014
rect 378520 335442 378548 338014
rect 378796 335782 378824 338014
rect 378784 335776 378836 335782
rect 378784 335718 378836 335724
rect 378508 335436 378560 335442
rect 378508 335378 378560 335384
rect 379072 335374 379100 338014
rect 379164 338014 379316 338042
rect 379592 338014 379744 338042
rect 379868 338014 380020 338042
rect 380144 338014 380388 338042
rect 378048 335368 378100 335374
rect 378048 335310 378100 335316
rect 379060 335368 379112 335374
rect 379060 335310 379112 335316
rect 377954 5128 378010 5137
rect 377954 5063 378010 5072
rect 378060 4894 378088 335310
rect 379164 7721 379192 338014
rect 379716 336161 379744 338014
rect 379702 336152 379758 336161
rect 379702 336087 379758 336096
rect 379992 335850 380020 338014
rect 380360 335918 380388 338014
rect 380498 337770 380526 338028
rect 380728 338014 380788 338042
rect 381064 338014 381216 338042
rect 381340 338014 381584 338042
rect 381708 338014 381860 338042
rect 381984 338014 382136 338042
rect 380498 337742 380572 337770
rect 380348 335912 380400 335918
rect 380348 335854 380400 335860
rect 379980 335844 380032 335850
rect 379980 335786 380032 335792
rect 379244 335776 379296 335782
rect 379296 335736 379468 335764
rect 379244 335718 379296 335724
rect 379244 335436 379296 335442
rect 379244 335378 379296 335384
rect 379150 7712 379206 7721
rect 379150 7647 379206 7656
rect 379256 6361 379284 335378
rect 379336 335368 379388 335374
rect 379336 335310 379388 335316
rect 379242 6352 379298 6361
rect 379242 6287 379298 6296
rect 377680 4888 377732 4894
rect 377680 4830 377732 4836
rect 378048 4888 378100 4894
rect 378048 4830 378100 4836
rect 376484 4072 376536 4078
rect 376484 4014 376536 4020
rect 375300 3590 375420 3618
rect 375196 3528 375248 3534
rect 375196 3470 375248 3476
rect 375392 3466 375420 3590
rect 375288 3460 375340 3466
rect 375288 3402 375340 3408
rect 375380 3460 375432 3466
rect 375380 3402 375432 3408
rect 375300 480 375328 3402
rect 376496 480 376524 4014
rect 377692 480 377720 4830
rect 379348 4826 379376 335310
rect 378876 4820 378928 4826
rect 378876 4762 378928 4768
rect 379336 4820 379388 4826
rect 379336 4762 379388 4768
rect 378888 480 378916 4762
rect 379440 3505 379468 335736
rect 380544 11830 380572 337742
rect 380624 335912 380676 335918
rect 380624 335854 380676 335860
rect 380532 11824 380584 11830
rect 380532 11766 380584 11772
rect 380636 7585 380664 335854
rect 380622 7576 380678 7585
rect 380622 7511 380678 7520
rect 380728 4865 380756 338014
rect 381188 335918 381216 338014
rect 381556 336297 381584 338014
rect 381542 336288 381598 336297
rect 381542 336223 381598 336232
rect 381176 335912 381228 335918
rect 381176 335854 381228 335860
rect 380808 335844 380860 335850
rect 380808 335786 380860 335792
rect 380820 5001 380848 335786
rect 381832 335354 381860 338014
rect 382108 336025 382136 338014
rect 382200 338014 382260 338042
rect 382094 336016 382150 336025
rect 382094 335951 382150 335960
rect 382096 335912 382148 335918
rect 382096 335854 382148 335860
rect 381832 335326 382044 335354
rect 382016 11762 382044 335326
rect 382004 11756 382056 11762
rect 382004 11698 382056 11704
rect 382108 6225 382136 335854
rect 382094 6216 382150 6225
rect 382094 6151 382150 6160
rect 380806 4992 380862 5001
rect 380806 4927 380862 4936
rect 380714 4856 380770 4865
rect 380714 4791 380770 4800
rect 381176 4208 381228 4214
rect 381176 4150 381228 4156
rect 379980 4004 380032 4010
rect 379980 3946 380032 3952
rect 379426 3496 379482 3505
rect 379426 3431 379482 3440
rect 379992 480 380020 3946
rect 381188 480 381216 4150
rect 382200 3369 382228 338014
rect 382936 46918 382964 487834
rect 383028 86970 383056 487970
rect 383120 126954 383148 488106
rect 383212 458182 383240 488378
rect 383384 488232 383436 488238
rect 383384 488174 383436 488180
rect 383292 486736 383344 486742
rect 383292 486678 383344 486684
rect 383200 458176 383252 458182
rect 383200 458118 383252 458124
rect 383200 335844 383252 335850
rect 383200 335786 383252 335792
rect 383108 126948 383160 126954
rect 383108 126890 383160 126896
rect 383016 86964 383068 86970
rect 383016 86906 383068 86912
rect 382924 46912 382976 46918
rect 382924 46854 382976 46860
rect 382372 6860 382424 6866
rect 382372 6802 382424 6808
rect 382186 3360 382242 3369
rect 382186 3295 382242 3304
rect 382384 480 382412 6802
rect 383212 2922 383240 335786
rect 383304 167006 383332 486678
rect 383396 206990 383424 488174
rect 383568 487008 383620 487014
rect 383568 486950 383620 486956
rect 383476 486940 383528 486946
rect 383476 486882 383528 486888
rect 383488 245614 383516 486882
rect 383580 299470 383608 486950
rect 384132 485790 384160 488446
rect 384212 487144 384264 487150
rect 384212 487086 384264 487092
rect 384120 485784 384172 485790
rect 384120 485726 384172 485732
rect 384224 405686 384252 487086
rect 384212 405680 384264 405686
rect 384212 405622 384264 405628
rect 383568 299464 383620 299470
rect 383568 299406 383620 299412
rect 383476 245608 383528 245614
rect 383476 245550 383528 245556
rect 383384 206984 383436 206990
rect 383384 206926 383436 206932
rect 383292 167000 383344 167006
rect 383292 166942 383344 166948
rect 384316 20670 384344 490039
rect 384486 489968 384542 489977
rect 384486 489903 384542 489912
rect 384396 486600 384448 486606
rect 384396 486542 384448 486548
rect 384408 73166 384436 486542
rect 384396 73160 384448 73166
rect 384396 73102 384448 73108
rect 384500 33114 384528 489903
rect 384672 488096 384724 488102
rect 384672 488038 384724 488044
rect 384580 487960 384632 487966
rect 384580 487902 384632 487908
rect 384592 113150 384620 487902
rect 384684 153202 384712 488038
rect 384948 487076 385000 487082
rect 384948 487018 385000 487024
rect 384856 486804 384908 486810
rect 384856 486746 384908 486752
rect 384764 486668 384816 486674
rect 384764 486610 384816 486616
rect 384776 193186 384804 486610
rect 384868 233238 384896 486746
rect 384960 353258 384988 487018
rect 384948 353252 385000 353258
rect 384948 353194 385000 353200
rect 384856 233232 384908 233238
rect 384856 233174 384908 233180
rect 384764 193180 384816 193186
rect 384764 193122 384816 193128
rect 384672 153196 384724 153202
rect 384672 153138 384724 153144
rect 384580 113144 384632 113150
rect 384580 113086 384632 113092
rect 385696 60722 385724 490175
rect 385868 488300 385920 488306
rect 385868 488242 385920 488248
rect 385776 486872 385828 486878
rect 385776 486814 385828 486820
rect 385788 273222 385816 486814
rect 385880 379506 385908 488242
rect 385972 419490 386000 490962
rect 386052 490952 386104 490958
rect 386052 490894 386104 490900
rect 386064 431934 386092 490894
rect 386144 488368 386196 488374
rect 386144 488310 386196 488316
rect 386156 471986 386184 488310
rect 393964 487824 394016 487830
rect 393964 487766 394016 487772
rect 386144 471980 386196 471986
rect 386144 471922 386196 471928
rect 386052 431928 386104 431934
rect 386052 431870 386104 431876
rect 385960 419484 386012 419490
rect 385960 419426 386012 419432
rect 385868 379500 385920 379506
rect 385868 379442 385920 379448
rect 391204 335980 391256 335986
rect 391204 335922 391256 335928
rect 385776 273216 385828 273222
rect 385776 273158 385828 273164
rect 385684 60716 385736 60722
rect 385684 60658 385736 60664
rect 384488 33108 384540 33114
rect 384488 33050 384540 33056
rect 384304 20664 384356 20670
rect 384304 20606 384356 20612
rect 391112 9920 391164 9926
rect 391112 9862 391164 9868
rect 389456 9852 389508 9858
rect 389456 9794 389508 9800
rect 387800 9784 387852 9790
rect 387800 9726 387852 9732
rect 384304 9716 384356 9722
rect 384304 9658 384356 9664
rect 383568 3936 383620 3942
rect 383568 3878 383620 3884
rect 383200 2916 383252 2922
rect 383200 2858 383252 2864
rect 383580 480 383608 3878
rect 384316 490 384344 9658
rect 385960 6996 386012 7002
rect 385960 6938 386012 6944
rect 384592 598 384804 626
rect 384592 490 384620 598
rect 335054 -960 335166 480
rect 336250 -960 336362 480
rect 337446 -960 337558 480
rect 338642 -960 338754 480
rect 339838 -960 339950 480
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 343334 -960 343446 480
rect 344530 -960 344642 480
rect 345726 -960 345838 480
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351614 -960 351726 480
rect 352810 -960 352922 480
rect 354006 -960 354118 480
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359894 -960 360006 480
rect 361090 -960 361202 480
rect 362286 -960 362398 480
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 368174 -960 368286 480
rect 369370 -960 369482 480
rect 370566 -960 370678 480
rect 371670 -960 371782 480
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376454 -960 376566 480
rect 377650 -960 377762 480
rect 378846 -960 378958 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384316 462 384620 490
rect 384776 480 384804 598
rect 385972 480 386000 6938
rect 387156 3868 387208 3874
rect 387156 3810 387208 3816
rect 387168 480 387196 3810
rect 387812 490 387840 9726
rect 388088 598 388300 626
rect 388088 490 388116 598
rect 384734 -960 384846 480
rect 385930 -960 386042 480
rect 387126 -960 387238 480
rect 387812 462 388116 490
rect 388272 480 388300 598
rect 389468 480 389496 9794
rect 390652 3732 390704 3738
rect 390652 3674 390704 3680
rect 390664 480 390692 3674
rect 391124 3482 391152 9862
rect 391216 3738 391244 335922
rect 392584 9988 392636 9994
rect 392584 9930 392636 9936
rect 391204 3732 391256 3738
rect 391204 3674 391256 3680
rect 391124 3454 391888 3482
rect 391860 480 391888 3454
rect 392596 490 392624 9930
rect 393976 6866 394004 487766
rect 580908 487756 580960 487762
rect 580908 487698 580960 487704
rect 580356 487688 580408 487694
rect 580356 487630 580408 487636
rect 580264 486192 580316 486198
rect 580264 486134 580316 486140
rect 580172 485784 580224 485790
rect 580172 485726 580224 485732
rect 580184 484673 580212 485726
rect 580170 484664 580226 484673
rect 580170 484599 580226 484608
rect 580172 471980 580224 471986
rect 580172 471922 580224 471928
rect 580184 471481 580212 471922
rect 580170 471472 580226 471481
rect 580170 471407 580226 471416
rect 580172 458176 580224 458182
rect 580170 458144 580172 458153
rect 580224 458144 580226 458153
rect 580170 458079 580226 458088
rect 580172 431928 580224 431934
rect 580172 431870 580224 431876
rect 580184 431633 580212 431870
rect 580170 431624 580226 431633
rect 580170 431559 580226 431568
rect 580172 419484 580224 419490
rect 580172 419426 580224 419432
rect 580184 418305 580212 419426
rect 580170 418296 580226 418305
rect 580170 418231 580226 418240
rect 580172 405680 580224 405686
rect 580172 405622 580224 405628
rect 580184 404977 580212 405622
rect 580170 404968 580226 404977
rect 580170 404903 580226 404912
rect 579988 379500 580040 379506
rect 579988 379442 580040 379448
rect 580000 378457 580028 379442
rect 579986 378448 580042 378457
rect 579986 378383 580042 378392
rect 580172 353252 580224 353258
rect 580172 353194 580224 353200
rect 580184 351937 580212 353194
rect 580170 351928 580226 351937
rect 580170 351863 580226 351872
rect 405096 336728 405148 336734
rect 405096 336670 405148 336676
rect 405004 335708 405056 335714
rect 405004 335650 405056 335656
rect 398104 335640 398156 335646
rect 398104 335582 398156 335588
rect 396724 335436 396776 335442
rect 396724 335378 396776 335384
rect 395344 10056 395396 10062
rect 395344 9998 395396 10004
rect 393964 6860 394016 6866
rect 393964 6802 394016 6808
rect 394238 4040 394294 4049
rect 394238 3975 394294 3984
rect 392872 598 393084 626
rect 392872 490 392900 598
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 392596 462 392900 490
rect 393056 480 393084 598
rect 394252 480 394280 3975
rect 395356 480 395384 9998
rect 396540 8356 396592 8362
rect 396540 8298 396592 8304
rect 396552 480 396580 8298
rect 396736 4146 396764 335378
rect 396724 4140 396776 4146
rect 396724 4082 396776 4088
rect 397734 3904 397790 3913
rect 397734 3839 397790 3848
rect 397748 480 397776 3839
rect 398116 3330 398144 335582
rect 403624 335572 403676 335578
rect 403624 335514 403676 335520
rect 399484 335504 399536 335510
rect 399484 335446 399536 335452
rect 398932 5568 398984 5574
rect 398932 5510 398984 5516
rect 398104 3324 398156 3330
rect 398104 3266 398156 3272
rect 398944 480 398972 5510
rect 399496 4078 399524 335446
rect 403532 8492 403584 8498
rect 403532 8434 403584 8440
rect 400128 8424 400180 8430
rect 400128 8366 400180 8372
rect 399484 4072 399536 4078
rect 399484 4014 399536 4020
rect 400140 480 400168 8366
rect 402520 5636 402572 5642
rect 402520 5578 402572 5584
rect 401322 3768 401378 3777
rect 401322 3703 401378 3712
rect 401336 480 401364 3703
rect 402532 480 402560 5578
rect 403544 3482 403572 8434
rect 403636 3942 403664 335514
rect 405016 4010 405044 335650
rect 405004 4004 405056 4010
rect 405004 3946 405056 3952
rect 403624 3936 403676 3942
rect 403624 3878 403676 3884
rect 404820 3664 404872 3670
rect 404820 3606 404872 3612
rect 403544 3454 403664 3482
rect 403636 480 403664 3454
rect 404832 480 404860 3606
rect 405108 2854 405136 336670
rect 417424 336660 417476 336666
rect 417424 336602 417476 336608
rect 416044 336524 416096 336530
rect 416044 336466 416096 336472
rect 411904 335844 411956 335850
rect 411904 335786 411956 335792
rect 410800 8628 410852 8634
rect 410800 8570 410852 8576
rect 407212 8560 407264 8566
rect 407212 8502 407264 8508
rect 406016 5704 406068 5710
rect 406016 5646 406068 5652
rect 405096 2848 405148 2854
rect 405096 2790 405148 2796
rect 406028 480 406056 5646
rect 407224 480 407252 8502
rect 409604 5772 409656 5778
rect 409604 5714 409656 5720
rect 408408 2916 408460 2922
rect 408408 2858 408460 2864
rect 408420 480 408448 2858
rect 409616 480 409644 5714
rect 410812 480 410840 8570
rect 411916 3874 411944 335786
rect 413284 335776 413336 335782
rect 413284 335718 413336 335724
rect 413100 5840 413152 5846
rect 413100 5782 413152 5788
rect 411904 3868 411956 3874
rect 411904 3810 411956 3816
rect 411902 3632 411958 3641
rect 411902 3567 411958 3576
rect 411916 480 411944 3567
rect 413112 480 413140 5782
rect 413296 3670 413324 335718
rect 414296 8696 414348 8702
rect 414296 8638 414348 8644
rect 413284 3664 413336 3670
rect 413284 3606 413336 3612
rect 414308 480 414336 8638
rect 416056 3738 416084 336466
rect 416688 5908 416740 5914
rect 416688 5850 416740 5856
rect 415492 3732 415544 3738
rect 415492 3674 415544 3680
rect 416044 3732 416096 3738
rect 416044 3674 416096 3680
rect 415504 480 415532 3674
rect 416700 480 416728 5850
rect 417436 2922 417464 336602
rect 425704 336592 425756 336598
rect 425704 336534 425756 336540
rect 418802 336424 418858 336433
rect 418802 336359 418858 336368
rect 417884 8764 417936 8770
rect 417884 8706 417936 8712
rect 417424 2916 417476 2922
rect 417424 2858 417476 2864
rect 417896 480 417924 8706
rect 418816 2922 418844 336359
rect 422942 336288 422998 336297
rect 422942 336223 422998 336232
rect 421380 8832 421432 8838
rect 421380 8774 421432 8780
rect 420184 5976 420236 5982
rect 420184 5918 420236 5924
rect 418804 2916 418856 2922
rect 418804 2858 418856 2864
rect 418620 2848 418672 2854
rect 418620 2790 418672 2796
rect 418632 490 418660 2790
rect 418816 598 419028 626
rect 418816 490 418844 598
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396510 -960 396622 480
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404790 -960 404902 480
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409574 -960 409686 480
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 413070 -960 413182 480
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417854 -960 417966 480
rect 418632 462 418844 490
rect 419000 480 419028 598
rect 420196 480 420224 5918
rect 421392 480 421420 8774
rect 422576 3732 422628 3738
rect 422576 3674 422628 3680
rect 422588 480 422616 3674
rect 422956 3641 422984 336223
rect 424968 8900 425020 8906
rect 424968 8842 425020 8848
rect 423772 6044 423824 6050
rect 423772 5986 423824 5992
rect 422942 3632 422998 3641
rect 422942 3567 422998 3576
rect 423784 480 423812 5986
rect 424980 480 425008 8842
rect 425716 3738 425744 336534
rect 429844 336456 429896 336462
rect 429844 336398 429896 336404
rect 425794 336152 425850 336161
rect 425794 336087 425850 336096
rect 425704 3732 425756 3738
rect 425704 3674 425756 3680
rect 425808 2786 425836 336087
rect 428464 9648 428516 9654
rect 428464 9590 428516 9596
rect 427268 6112 427320 6118
rect 427268 6054 427320 6060
rect 426164 3800 426216 3806
rect 426164 3742 426216 3748
rect 425796 2780 425848 2786
rect 425796 2722 425848 2728
rect 426176 480 426204 3742
rect 427280 480 427308 6054
rect 428476 480 428504 9590
rect 429856 3806 429884 336398
rect 432604 336388 432656 336394
rect 432604 336330 432656 336336
rect 432052 9580 432104 9586
rect 432052 9522 432104 9528
rect 430856 6792 430908 6798
rect 430856 6734 430908 6740
rect 429844 3800 429896 3806
rect 429844 3742 429896 3748
rect 429660 2984 429712 2990
rect 429660 2926 429712 2932
rect 429672 480 429700 2926
rect 430868 480 430896 6734
rect 432064 480 432092 9522
rect 432616 3806 432644 336330
rect 436744 336320 436796 336326
rect 436744 336262 436796 336268
rect 436756 16574 436784 336262
rect 440884 336252 440936 336258
rect 440884 336194 440936 336200
rect 436756 16546 436968 16574
rect 435548 9512 435600 9518
rect 435548 9454 435600 9460
rect 434444 6724 434496 6730
rect 434444 6666 434496 6672
rect 432512 3800 432564 3806
rect 432512 3742 432564 3748
rect 432604 3800 432656 3806
rect 432604 3742 432656 3748
rect 432524 2922 432552 3742
rect 432512 2916 432564 2922
rect 432512 2858 432564 2864
rect 433248 2916 433300 2922
rect 433248 2858 433300 2864
rect 433260 480 433288 2858
rect 434456 480 434484 6666
rect 435560 480 435588 9454
rect 436744 3052 436796 3058
rect 436744 2994 436796 3000
rect 436756 480 436784 2994
rect 436940 2990 436968 16546
rect 439136 9444 439188 9450
rect 439136 9386 439188 9392
rect 437940 6656 437992 6662
rect 437940 6598 437992 6604
rect 436928 2984 436980 2990
rect 436928 2926 436980 2932
rect 437952 480 437980 6598
rect 439148 480 439176 9386
rect 440332 3800 440384 3806
rect 440332 3742 440384 3748
rect 440344 480 440372 3742
rect 440896 3058 440924 336194
rect 443644 336184 443696 336190
rect 443644 336126 443696 336132
rect 443656 16574 443684 336126
rect 447784 336116 447836 336122
rect 447784 336058 447836 336064
rect 443656 16546 443960 16574
rect 442632 9376 442684 9382
rect 442632 9318 442684 9324
rect 441528 6588 441580 6594
rect 441528 6530 441580 6536
rect 440884 3052 440936 3058
rect 440884 2994 440936 3000
rect 441540 480 441568 6530
rect 442644 480 442672 9318
rect 443932 3126 443960 16546
rect 446220 9308 446272 9314
rect 446220 9250 446272 9256
rect 445024 6520 445076 6526
rect 445024 6462 445076 6468
rect 443828 3120 443880 3126
rect 443828 3062 443880 3068
rect 443920 3120 443972 3126
rect 443920 3062 443972 3068
rect 443840 480 443868 3062
rect 445036 480 445064 6462
rect 446232 480 446260 9250
rect 447796 3058 447824 336058
rect 450544 336048 450596 336054
rect 450544 335990 450596 335996
rect 451922 336016 451978 336025
rect 450556 16574 450584 335990
rect 451922 335951 451978 335960
rect 450556 16546 451044 16574
rect 449808 9240 449860 9246
rect 449808 9182 449860 9188
rect 448612 6452 448664 6458
rect 448612 6394 448664 6400
rect 447784 3052 447836 3058
rect 447784 2994 447836 3000
rect 447416 2984 447468 2990
rect 447416 2926 447468 2932
rect 447428 480 447456 2926
rect 448624 480 448652 6394
rect 449820 480 449848 9182
rect 451016 2854 451044 16546
rect 451936 3777 451964 335951
rect 580172 299464 580224 299470
rect 580172 299406 580224 299412
rect 580184 298761 580212 299406
rect 580170 298752 580226 298761
rect 580170 298687 580226 298696
rect 580172 273216 580224 273222
rect 580172 273158 580224 273164
rect 580184 272241 580212 273158
rect 580170 272232 580226 272241
rect 580170 272167 580226 272176
rect 580172 245608 580224 245614
rect 580170 245576 580172 245585
rect 580224 245576 580226 245585
rect 580170 245511 580226 245520
rect 579988 233232 580040 233238
rect 579988 233174 580040 233180
rect 580000 232393 580028 233174
rect 579986 232384 580042 232393
rect 579986 232319 580042 232328
rect 580172 206984 580224 206990
rect 580172 206926 580224 206932
rect 580184 205737 580212 206926
rect 580170 205728 580226 205737
rect 580170 205663 580226 205672
rect 580172 193180 580224 193186
rect 580172 193122 580224 193128
rect 580184 192545 580212 193122
rect 580170 192536 580226 192545
rect 580170 192471 580226 192480
rect 580172 167000 580224 167006
rect 580172 166942 580224 166948
rect 580184 165889 580212 166942
rect 580170 165880 580226 165889
rect 580170 165815 580226 165824
rect 579620 153196 579672 153202
rect 579620 153138 579672 153144
rect 579632 152697 579660 153138
rect 579618 152688 579674 152697
rect 579618 152623 579674 152632
rect 580172 126948 580224 126954
rect 580172 126890 580224 126896
rect 580184 126041 580212 126890
rect 580170 126032 580226 126041
rect 580170 125967 580226 125976
rect 580172 113144 580224 113150
rect 580172 113086 580224 113092
rect 580184 112849 580212 113086
rect 580170 112840 580226 112849
rect 580170 112775 580226 112784
rect 580276 99521 580304 486134
rect 580368 139369 580396 487630
rect 580724 486532 580776 486538
rect 580724 486474 580776 486480
rect 580632 486396 580684 486402
rect 580632 486338 580684 486344
rect 580540 486328 580592 486334
rect 580540 486270 580592 486276
rect 580448 486260 580500 486266
rect 580448 486202 580500 486208
rect 580460 179217 580488 486202
rect 580552 219065 580580 486270
rect 580644 258913 580672 486338
rect 580736 312089 580764 486474
rect 580816 486464 580868 486470
rect 580816 486406 580868 486412
rect 580828 325281 580856 486406
rect 580920 365129 580948 487698
rect 580906 365120 580962 365129
rect 580906 365055 580962 365064
rect 580814 325272 580870 325281
rect 580814 325207 580870 325216
rect 580722 312080 580778 312089
rect 580722 312015 580778 312024
rect 580630 258904 580686 258913
rect 580630 258839 580686 258848
rect 580538 219056 580594 219065
rect 580538 218991 580594 219000
rect 580446 179208 580502 179217
rect 580446 179143 580502 179152
rect 580354 139360 580410 139369
rect 580354 139295 580410 139304
rect 580262 99512 580318 99521
rect 580262 99447 580318 99456
rect 580172 86964 580224 86970
rect 580172 86906 580224 86912
rect 580184 86193 580212 86906
rect 580170 86184 580226 86193
rect 580170 86119 580226 86128
rect 580172 73160 580224 73166
rect 580172 73102 580224 73108
rect 580184 73001 580212 73102
rect 580170 72992 580226 73001
rect 580170 72927 580226 72936
rect 580172 60716 580224 60722
rect 580172 60658 580224 60664
rect 580184 59673 580212 60658
rect 580170 59664 580226 59673
rect 580170 59599 580226 59608
rect 580172 46912 580224 46918
rect 580172 46854 580224 46860
rect 580184 46345 580212 46854
rect 580170 46336 580226 46345
rect 580170 46271 580226 46280
rect 580170 33144 580226 33153
rect 580170 33079 580172 33088
rect 580224 33079 580226 33088
rect 580172 33050 580224 33056
rect 579988 20664 580040 20670
rect 579988 20606 580040 20612
rect 580000 19825 580028 20606
rect 579986 19816 580042 19825
rect 579986 19751 580042 19760
rect 503720 12232 503772 12238
rect 503720 12174 503772 12180
rect 480536 11008 480588 11014
rect 480536 10950 480588 10956
rect 476488 10260 476540 10266
rect 476488 10202 476540 10208
rect 473452 10192 473504 10198
rect 473452 10134 473504 10140
rect 473360 10124 473412 10130
rect 473360 10066 473412 10072
rect 467470 9208 467526 9217
rect 453304 9172 453356 9178
rect 467470 9143 467526 9152
rect 453304 9114 453356 9120
rect 452108 6384 452160 6390
rect 452108 6326 452160 6332
rect 451922 3768 451978 3777
rect 451922 3703 451978 3712
rect 450912 2848 450964 2854
rect 450912 2790 450964 2796
rect 451004 2848 451056 2854
rect 451004 2790 451056 2796
rect 450924 480 450952 2790
rect 452120 480 452148 6326
rect 453316 480 453344 9114
rect 456892 9104 456944 9110
rect 456892 9046 456944 9052
rect 455696 6316 455748 6322
rect 455696 6258 455748 6264
rect 454500 3120 454552 3126
rect 454500 3062 454552 3068
rect 454512 480 454540 3062
rect 455708 480 455736 6258
rect 456904 480 456932 9046
rect 460388 9036 460440 9042
rect 460388 8978 460440 8984
rect 459192 6248 459244 6254
rect 459192 6190 459244 6196
rect 458088 3188 458140 3194
rect 458088 3130 458140 3136
rect 458100 480 458128 3130
rect 459204 480 459232 6190
rect 460400 480 460428 8978
rect 463976 8968 464028 8974
rect 463976 8910 464028 8916
rect 462780 6180 462832 6186
rect 462780 6122 462832 6128
rect 461584 2984 461636 2990
rect 461584 2926 461636 2932
rect 461596 480 461624 2926
rect 462792 480 462820 6122
rect 463988 480 464016 8910
rect 466274 6624 466330 6633
rect 466274 6559 466330 6568
rect 465172 3256 465224 3262
rect 465172 3198 465224 3204
rect 465184 480 465212 3198
rect 466288 480 466316 6559
rect 467484 480 467512 9143
rect 471058 9072 471114 9081
rect 471058 9007 471114 9016
rect 469862 6488 469918 6497
rect 469862 6423 469918 6432
rect 468668 3052 468720 3058
rect 468668 2994 468720 3000
rect 468680 480 468708 2994
rect 469876 480 469904 6423
rect 471072 480 471100 9007
rect 473372 3398 473400 10066
rect 472256 3392 472308 3398
rect 472256 3334 472308 3340
rect 473360 3392 473412 3398
rect 473360 3334 473412 3340
rect 472268 480 472296 3334
rect 473464 480 473492 10134
rect 474556 3392 474608 3398
rect 474556 3334 474608 3340
rect 474568 480 474596 3334
rect 475752 2848 475804 2854
rect 475752 2790 475804 2796
rect 475764 480 475792 2790
rect 476500 490 476528 10202
rect 478142 8936 478198 8945
rect 478142 8871 478198 8880
rect 476776 598 476988 626
rect 476776 490 476804 598
rect 418958 -960 419070 480
rect 420154 -960 420266 480
rect 421350 -960 421462 480
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 426134 -960 426246 480
rect 427238 -960 427350 480
rect 428434 -960 428546 480
rect 429630 -960 429742 480
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 434414 -960 434526 480
rect 435518 -960 435630 480
rect 436714 -960 436826 480
rect 437910 -960 438022 480
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443798 -960 443910 480
rect 444994 -960 445106 480
rect 446190 -960 446302 480
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 452078 -960 452190 480
rect 453274 -960 453386 480
rect 454470 -960 454582 480
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 460358 -960 460470 480
rect 461554 -960 461666 480
rect 462750 -960 462862 480
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 466246 -960 466358 480
rect 467442 -960 467554 480
rect 468638 -960 468750 480
rect 469834 -960 469946 480
rect 471030 -960 471142 480
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474526 -960 474638 480
rect 475722 -960 475834 480
rect 476500 462 476804 490
rect 476960 480 476988 598
rect 478156 480 478184 8871
rect 479340 2916 479392 2922
rect 479340 2858 479392 2864
rect 479352 480 479380 2858
rect 480548 480 480576 10950
rect 481640 10940 481692 10946
rect 481640 10882 481692 10888
rect 481652 3398 481680 10882
rect 481732 10872 481784 10878
rect 481732 10814 481784 10820
rect 481640 3392 481692 3398
rect 481640 3334 481692 3340
rect 481744 480 481772 10814
rect 484768 10804 484820 10810
rect 484768 10746 484820 10752
rect 484032 10736 484084 10742
rect 484032 10678 484084 10684
rect 482836 3392 482888 3398
rect 482836 3334 482888 3340
rect 482848 480 482876 3334
rect 484044 480 484072 10678
rect 484780 490 484808 10746
rect 486424 10668 486476 10674
rect 486424 10610 486476 10616
rect 485056 598 485268 626
rect 485056 490 485084 598
rect 476918 -960 477030 480
rect 478114 -960 478226 480
rect 479310 -960 479422 480
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482806 -960 482918 480
rect 484002 -960 484114 480
rect 484780 462 485084 490
rect 485240 480 485268 598
rect 486436 480 486464 10610
rect 487160 10600 487212 10606
rect 487160 10542 487212 10548
rect 494702 10568 494758 10577
rect 487172 490 487200 10542
rect 488816 10532 488868 10538
rect 494702 10503 494758 10512
rect 488816 10474 488868 10480
rect 487448 598 487660 626
rect 487448 490 487476 598
rect 485198 -960 485310 480
rect 486394 -960 486506 480
rect 487172 462 487476 490
rect 487632 480 487660 598
rect 488828 480 488856 10474
rect 490012 10464 490064 10470
rect 490012 10406 490064 10412
rect 489920 10396 489972 10402
rect 489920 10338 489972 10344
rect 489932 4214 489960 10338
rect 489920 4208 489972 4214
rect 489920 4150 489972 4156
rect 490024 3482 490052 10406
rect 493048 10328 493100 10334
rect 493048 10270 493100 10276
rect 492312 7064 492364 7070
rect 492312 7006 492364 7012
rect 491116 4208 491168 4214
rect 491116 4150 491168 4156
rect 489932 3454 490052 3482
rect 489932 480 489960 3454
rect 491128 480 491156 4150
rect 492324 480 492352 7006
rect 493060 490 493088 10270
rect 493336 598 493548 626
rect 493336 490 493364 598
rect 487590 -960 487702 480
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 491086 -960 491198 480
rect 492282 -960 492394 480
rect 493060 462 493364 490
rect 493520 480 493548 598
rect 494716 480 494744 10503
rect 497094 10432 497150 10441
rect 497094 10367 497150 10376
rect 495900 7132 495952 7138
rect 495900 7074 495952 7080
rect 495912 480 495940 7074
rect 497108 480 497136 10367
rect 500590 10296 500646 10305
rect 500590 10231 500646 10240
rect 499396 7200 499448 7206
rect 499396 7142 499448 7148
rect 498200 4276 498252 4282
rect 498200 4218 498252 4224
rect 498212 480 498240 4218
rect 499408 480 499436 7142
rect 500604 480 500632 10231
rect 502984 7268 503036 7274
rect 502984 7210 503036 7216
rect 501788 4344 501840 4350
rect 501788 4286 501840 4292
rect 501800 480 501828 4286
rect 502996 480 503024 7210
rect 503732 490 503760 12174
rect 507216 12164 507268 12170
rect 507216 12106 507268 12112
rect 506480 7336 506532 7342
rect 506480 7278 506532 7284
rect 505376 4412 505428 4418
rect 505376 4354 505428 4360
rect 504008 598 504220 626
rect 504008 490 504036 598
rect 493478 -960 493590 480
rect 494674 -960 494786 480
rect 495870 -960 495982 480
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 499366 -960 499478 480
rect 500562 -960 500674 480
rect 501758 -960 501870 480
rect 502954 -960 503066 480
rect 503732 462 504036 490
rect 504192 480 504220 598
rect 505388 480 505416 4354
rect 506492 480 506520 7278
rect 507228 490 507256 12106
rect 517888 12096 517940 12102
rect 517888 12038 517940 12044
rect 511262 10704 511318 10713
rect 511262 10639 511318 10648
rect 510068 7404 510120 7410
rect 510068 7346 510120 7352
rect 508872 4480 508924 4486
rect 508872 4422 508924 4428
rect 507504 598 507716 626
rect 507504 490 507532 598
rect 504150 -960 504262 480
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507228 462 507532 490
rect 507688 480 507716 598
rect 508884 480 508912 4422
rect 510080 480 510108 7346
rect 511276 480 511304 10639
rect 517152 7540 517204 7546
rect 517152 7482 517204 7488
rect 513564 7472 513616 7478
rect 513564 7414 513616 7420
rect 512460 4548 512512 4554
rect 512460 4490 512512 4496
rect 512472 480 512500 4490
rect 513576 480 513604 7414
rect 515956 4616 516008 4622
rect 515956 4558 516008 4564
rect 514760 3324 514812 3330
rect 514760 3266 514812 3272
rect 514772 480 514800 3266
rect 515968 480 515996 4558
rect 517164 480 517192 7482
rect 517900 490 517928 12038
rect 525432 12028 525484 12034
rect 525432 11970 525484 11976
rect 520740 8288 520792 8294
rect 520740 8230 520792 8236
rect 519544 4684 519596 4690
rect 519544 4626 519596 4632
rect 518176 598 518388 626
rect 518176 490 518204 598
rect 507646 -960 507758 480
rect 508842 -960 508954 480
rect 510038 -960 510150 480
rect 511234 -960 511346 480
rect 512430 -960 512542 480
rect 513534 -960 513646 480
rect 514730 -960 514842 480
rect 515926 -960 516038 480
rect 517122 -960 517234 480
rect 517900 462 518204 490
rect 518360 480 518388 598
rect 519556 480 519584 4626
rect 520752 480 520780 8230
rect 524236 8220 524288 8226
rect 524236 8162 524288 8168
rect 523040 4752 523092 4758
rect 523040 4694 523092 4700
rect 521844 4140 521896 4146
rect 521844 4082 521896 4088
rect 521856 480 521884 4082
rect 523052 480 523080 4694
rect 524248 480 524276 8162
rect 525444 480 525472 11970
rect 539600 11960 539652 11966
rect 539600 11902 539652 11908
rect 527824 8152 527876 8158
rect 527824 8094 527876 8100
rect 526628 5500 526680 5506
rect 526628 5442 526680 5448
rect 526640 480 526668 5442
rect 527836 480 527864 8094
rect 531320 8084 531372 8090
rect 531320 8026 531372 8032
rect 530124 5432 530176 5438
rect 530124 5374 530176 5380
rect 529020 4072 529072 4078
rect 529020 4014 529072 4020
rect 529032 480 529060 4014
rect 530136 480 530164 5374
rect 531332 480 531360 8026
rect 534908 8016 534960 8022
rect 534908 7958 534960 7964
rect 533712 5364 533764 5370
rect 533712 5306 533764 5312
rect 532516 3596 532568 3602
rect 532516 3538 532568 3544
rect 532528 480 532556 3538
rect 533724 480 533752 5306
rect 534920 480 534948 7958
rect 538404 7948 538456 7954
rect 538404 7890 538456 7896
rect 537208 5296 537260 5302
rect 537208 5238 537260 5244
rect 536104 4004 536156 4010
rect 536104 3946 536156 3952
rect 536116 480 536144 3946
rect 537220 480 537248 5238
rect 538416 480 538444 7890
rect 539612 480 539640 11902
rect 546684 11892 546736 11898
rect 546684 11834 546736 11840
rect 541992 7880 542044 7886
rect 541992 7822 542044 7828
rect 540796 5228 540848 5234
rect 540796 5170 540848 5176
rect 540808 480 540836 5170
rect 542004 480 542032 7822
rect 545488 7812 545540 7818
rect 545488 7754 545540 7760
rect 544384 5160 544436 5166
rect 544384 5102 544436 5108
rect 543188 3936 543240 3942
rect 543188 3878 543240 3884
rect 543200 480 543228 3878
rect 544396 480 544424 5102
rect 545500 480 545528 7754
rect 546696 480 546724 11834
rect 575112 11824 575164 11830
rect 575112 11766 575164 11772
rect 559746 7984 559802 7993
rect 559746 7919 559802 7928
rect 549076 7744 549128 7750
rect 549076 7686 549128 7692
rect 547880 5092 547932 5098
rect 547880 5034 547932 5040
rect 547892 480 547920 5034
rect 549088 480 549116 7686
rect 552664 7676 552716 7682
rect 552664 7618 552716 7624
rect 551468 5024 551520 5030
rect 551468 4966 551520 4972
rect 550272 3528 550324 3534
rect 550272 3470 550324 3476
rect 550284 480 550312 3470
rect 551480 480 551508 4966
rect 552676 480 552704 7618
rect 556160 7608 556212 7614
rect 556160 7550 556212 7556
rect 554964 4956 555016 4962
rect 554964 4898 555016 4904
rect 553768 3460 553820 3466
rect 553768 3402 553820 3408
rect 553780 480 553808 3402
rect 554976 480 555004 4898
rect 556172 480 556200 7550
rect 558550 5264 558606 5273
rect 558550 5199 558606 5208
rect 557356 3868 557408 3874
rect 557356 3810 557408 3816
rect 557368 480 557396 3810
rect 558564 480 558592 5199
rect 559760 480 559788 7919
rect 563242 7848 563298 7857
rect 563242 7783 563298 7792
rect 562048 4888 562100 4894
rect 562048 4830 562100 4836
rect 560852 3664 560904 3670
rect 560852 3606 560904 3612
rect 560864 480 560892 3606
rect 562060 480 562088 4830
rect 563256 480 563284 7783
rect 570326 7712 570382 7721
rect 570326 7647 570382 7656
rect 566830 6352 566886 6361
rect 566830 6287 566886 6296
rect 565634 5128 565690 5137
rect 565634 5063 565690 5072
rect 564440 3732 564492 3738
rect 564440 3674 564492 3680
rect 564452 480 564480 3674
rect 565648 480 565676 5063
rect 566844 480 566872 6287
rect 569132 4820 569184 4826
rect 569132 4762 569184 4768
rect 568026 3496 568082 3505
rect 568026 3431 568082 3440
rect 568040 480 568068 3431
rect 569144 480 569172 4762
rect 570340 480 570368 7647
rect 573914 7576 573970 7585
rect 573914 7511 573970 7520
rect 572718 4992 572774 5001
rect 572718 4927 572774 4936
rect 571524 3800 571576 3806
rect 571524 3742 571576 3748
rect 571536 480 571564 3742
rect 572732 480 572760 4927
rect 573928 480 573956 7511
rect 575124 480 575152 11766
rect 581000 11756 581052 11762
rect 581000 11698 581052 11704
rect 580172 6860 580224 6866
rect 580172 6802 580224 6808
rect 580184 6633 580212 6802
rect 580170 6624 580226 6633
rect 580170 6559 580226 6568
rect 577410 6216 577466 6225
rect 577410 6151 577466 6160
rect 576306 4856 576362 4865
rect 576306 4791 576362 4800
rect 576320 480 576348 4791
rect 577424 480 577452 6151
rect 578606 3632 578662 3641
rect 578606 3567 578662 3576
rect 578620 480 578648 3567
rect 581012 480 581040 11698
rect 582194 3768 582250 3777
rect 582194 3703 582250 3712
rect 582208 480 582236 3703
rect 583390 3360 583446 3369
rect 583390 3295 583446 3304
rect 583404 480 583432 3295
rect 518318 -960 518430 480
rect 519514 -960 519626 480
rect 520710 -960 520822 480
rect 521814 -960 521926 480
rect 523010 -960 523122 480
rect 524206 -960 524318 480
rect 525402 -960 525514 480
rect 526598 -960 526710 480
rect 527794 -960 527906 480
rect 528990 -960 529102 480
rect 530094 -960 530206 480
rect 531290 -960 531402 480
rect 532486 -960 532598 480
rect 533682 -960 533794 480
rect 534878 -960 534990 480
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538374 -960 538486 480
rect 539570 -960 539682 480
rect 540766 -960 540878 480
rect 541962 -960 542074 480
rect 543158 -960 543270 480
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546654 -960 546766 480
rect 547850 -960 547962 480
rect 549046 -960 549158 480
rect 550242 -960 550354 480
rect 551438 -960 551550 480
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554934 -960 555046 480
rect 556130 -960 556242 480
rect 557326 -960 557438 480
rect 558522 -960 558634 480
rect 559718 -960 559830 480
rect 560822 -960 560934 480
rect 562018 -960 562130 480
rect 563214 -960 563326 480
rect 564410 -960 564522 480
rect 565606 -960 565718 480
rect 566802 -960 566914 480
rect 567998 -960 568110 480
rect 569102 -960 569214 480
rect 570298 -960 570410 480
rect 571494 -960 571606 480
rect 572690 -960 572802 480
rect 573886 -960 573998 480
rect 575082 -960 575194 480
rect 576278 -960 576390 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 40498 700576 40554 700632
rect 24306 700440 24362 700496
rect 8114 700304 8170 700360
rect 3422 684256 3478 684312
rect 3514 671200 3570 671256
rect 3422 658144 3478 658200
rect 3422 632068 3424 632088
rect 3424 632068 3476 632088
rect 3476 632068 3478 632088
rect 3422 632032 3478 632068
rect 3146 619112 3202 619168
rect 3238 606056 3294 606112
rect 3330 579944 3386 580000
rect 3422 566888 3478 566944
rect 3422 553832 3478 553888
rect 3422 527856 3478 527912
rect 3422 514820 3478 514856
rect 3422 514800 3424 514820
rect 3424 514800 3476 514820
rect 3476 514800 3478 514820
rect 3054 501744 3110 501800
rect 2778 475668 2780 475688
rect 2780 475668 2832 475688
rect 2832 475668 2834 475688
rect 2778 475632 2834 475668
rect 3238 462576 3294 462632
rect 3238 449556 3240 449576
rect 3240 449556 3292 449576
rect 3292 449556 3294 449576
rect 3238 449520 3294 449556
rect 2778 423580 2780 423600
rect 2780 423580 2832 423600
rect 2832 423580 2834 423600
rect 2778 423544 2834 423580
rect 3330 410488 3386 410544
rect 2778 397432 2834 397488
rect 2778 371320 2834 371376
rect 2778 319232 2834 319288
rect 3146 293120 3202 293176
rect 2778 267144 2834 267200
rect 3238 241068 3240 241088
rect 3240 241068 3292 241088
rect 3292 241068 3294 241088
rect 3238 241032 3294 241068
rect 3238 188844 3240 188864
rect 3240 188844 3292 188864
rect 3292 188844 3294 188864
rect 3238 188808 3294 188844
rect 4066 358400 4122 358456
rect 3974 345344 4030 345400
rect 3882 306176 3938 306232
rect 3790 254088 3846 254144
rect 3698 214920 3754 214976
rect 3606 201864 3662 201920
rect 3514 162832 3570 162888
rect 3422 149776 3478 149832
rect 3238 136720 3294 136776
rect 2778 110608 2834 110664
rect 3330 97552 3386 97608
rect 2778 84632 2834 84688
rect 2778 71612 2780 71632
rect 2780 71612 2832 71632
rect 2832 71612 2834 71632
rect 2778 71576 2834 71612
rect 3054 58520 3110 58576
rect 3422 45500 3424 45520
rect 3424 45500 3476 45520
rect 3476 45500 3478 45520
rect 3422 45464 3478 45500
rect 6182 485968 6238 486024
rect 5446 335960 5502 336016
rect 2778 32408 2834 32464
rect 3054 19352 3110 19408
rect 1306 11600 1362 11656
rect 3422 6432 3478 6488
rect 7838 485832 7894 485888
rect 242438 490184 242494 490240
rect 238574 490048 238630 490104
rect 237286 489912 237342 489968
rect 293866 700712 293922 700768
rect 324318 700576 324374 700632
rect 319442 700440 319498 700496
rect 325698 700304 325754 700360
rect 559654 700712 559710 700768
rect 580170 697176 580226 697232
rect 580170 683848 580226 683904
rect 580170 670656 580226 670712
rect 580170 644000 580226 644056
rect 580170 630808 580226 630864
rect 580170 617480 580226 617536
rect 579802 590960 579858 591016
rect 580170 577632 580226 577688
rect 579802 564304 579858 564360
rect 580170 537784 580226 537840
rect 580170 524476 580226 524512
rect 580170 524456 580172 524476
rect 580172 524456 580224 524476
rect 580224 524456 580226 524476
rect 580170 511264 580226 511320
rect 385682 490184 385738 490240
rect 384302 490048 384358 490104
rect 373906 487056 373962 487112
rect 372618 486920 372674 486976
rect 377586 486920 377642 486976
rect 8022 486104 8078 486160
rect 12346 336232 12402 336288
rect 10966 336096 11022 336152
rect 8758 7520 8814 7576
rect 6458 3304 6514 3360
rect 12254 7656 12310 7712
rect 13542 10240 13598 10296
rect 17038 7792 17094 7848
rect 14738 3576 14794 3632
rect 15934 3440 15990 3496
rect 19430 3712 19486 3768
rect 26514 8880 26570 8936
rect 21822 7928 21878 7984
rect 30102 9016 30158 9072
rect 37002 10376 37058 10432
rect 41326 10512 41382 10568
rect 45466 10648 45522 10704
rect 47858 6160 47914 6216
rect 51354 6296 51410 6352
rect 54942 6432 54998 6488
rect 58438 6568 58494 6624
rect 79690 12008 79746 12064
rect 78586 11736 78642 11792
rect 81346 11872 81402 11928
rect 135258 9288 135314 9344
rect 131762 9152 131818 9208
rect 129370 4800 129426 4856
rect 132958 4936 133014 4992
rect 168378 5208 168434 5264
rect 175462 5072 175518 5128
rect 234618 11600 234674 11656
rect 236090 335960 236146 336016
rect 237654 336232 237710 336288
rect 237378 336096 237434 336152
rect 236182 7520 236238 7576
rect 236274 3304 236330 3360
rect 237562 10240 237618 10296
rect 237470 7656 237526 7712
rect 237378 3576 237434 3632
rect 238942 7792 238998 7848
rect 238850 3712 238906 3768
rect 239034 3440 239090 3496
rect 240414 7928 240470 7984
rect 241794 9016 241850 9072
rect 241702 8880 241758 8936
rect 243542 5208 243598 5264
rect 240506 3440 240562 3496
rect 239310 3304 239366 3360
rect 244554 10512 244610 10568
rect 244462 10376 244518 10432
rect 245842 10648 245898 10704
rect 247222 6296 247278 6352
rect 247130 6160 247186 6216
rect 248510 6568 248566 6624
rect 248602 6432 248658 6488
rect 254122 12008 254178 12064
rect 254214 11736 254270 11792
rect 255502 11872 255558 11928
rect 260654 3576 260710 3632
rect 266726 4800 266782 4856
rect 268014 9152 268070 9208
rect 269302 9288 269358 9344
rect 267738 4936 267794 4992
rect 267738 3712 267794 3768
rect 278778 5072 278834 5128
rect 295430 3440 295486 3496
rect 295522 3304 295578 3360
rect 300950 3576 301006 3632
rect 302514 3712 302570 3768
rect 332230 330520 332286 330576
rect 332414 330520 332470 330576
rect 335266 3984 335322 4040
rect 336554 3848 336610 3904
rect 336646 3712 336702 3768
rect 339406 3576 339462 3632
rect 352930 9152 352986 9208
rect 353022 6568 353078 6624
rect 354402 9016 354458 9072
rect 354494 6432 354550 6488
rect 360014 10512 360070 10568
rect 355966 8880 356022 8936
rect 361210 10376 361266 10432
rect 362590 10240 362646 10296
rect 376574 7928 376630 7984
rect 377862 336368 377918 336424
rect 377402 10648 377458 10704
rect 377862 7792 377918 7848
rect 376666 5208 376722 5264
rect 377954 5072 378010 5128
rect 379702 336096 379758 336152
rect 379150 7656 379206 7712
rect 379242 6296 379298 6352
rect 380622 7520 380678 7576
rect 381542 336232 381598 336288
rect 382094 335960 382150 336016
rect 382094 6160 382150 6216
rect 380806 4936 380862 4992
rect 380714 4800 380770 4856
rect 379426 3440 379482 3496
rect 382186 3304 382242 3360
rect 384486 489912 384542 489968
rect 580170 484608 580226 484664
rect 580170 471416 580226 471472
rect 580170 458124 580172 458144
rect 580172 458124 580224 458144
rect 580224 458124 580226 458144
rect 580170 458088 580226 458124
rect 580170 431568 580226 431624
rect 580170 418240 580226 418296
rect 580170 404912 580226 404968
rect 579986 378392 580042 378448
rect 580170 351872 580226 351928
rect 394238 3984 394294 4040
rect 397734 3848 397790 3904
rect 401322 3712 401378 3768
rect 411902 3576 411958 3632
rect 418802 336368 418858 336424
rect 422942 336232 422998 336288
rect 422942 3576 422998 3632
rect 425794 336096 425850 336152
rect 451922 335960 451978 336016
rect 580170 298696 580226 298752
rect 580170 272176 580226 272232
rect 580170 245556 580172 245576
rect 580172 245556 580224 245576
rect 580224 245556 580226 245576
rect 580170 245520 580226 245556
rect 579986 232328 580042 232384
rect 580170 205672 580226 205728
rect 580170 192480 580226 192536
rect 580170 165824 580226 165880
rect 579618 152632 579674 152688
rect 580170 125976 580226 126032
rect 580170 112784 580226 112840
rect 580906 365064 580962 365120
rect 580814 325216 580870 325272
rect 580722 312024 580778 312080
rect 580630 258848 580686 258904
rect 580538 219000 580594 219056
rect 580446 179152 580502 179208
rect 580354 139304 580410 139360
rect 580262 99456 580318 99512
rect 580170 86128 580226 86184
rect 580170 72936 580226 72992
rect 580170 59608 580226 59664
rect 580170 46280 580226 46336
rect 580170 33108 580226 33144
rect 580170 33088 580172 33108
rect 580172 33088 580224 33108
rect 580224 33088 580226 33108
rect 579986 19760 580042 19816
rect 467470 9152 467526 9208
rect 451922 3712 451978 3768
rect 466274 6568 466330 6624
rect 471058 9016 471114 9072
rect 469862 6432 469918 6488
rect 478142 8880 478198 8936
rect 494702 10512 494758 10568
rect 497094 10376 497150 10432
rect 500590 10240 500646 10296
rect 511262 10648 511318 10704
rect 559746 7928 559802 7984
rect 558550 5208 558606 5264
rect 563242 7792 563298 7848
rect 570326 7656 570382 7712
rect 566830 6296 566886 6352
rect 565634 5072 565690 5128
rect 568026 3440 568082 3496
rect 573914 7520 573970 7576
rect 572718 4936 572774 4992
rect 580170 6568 580226 6624
rect 577410 6160 577466 6216
rect 576306 4800 576362 4856
rect 578606 3576 578662 3632
rect 582194 3712 582250 3768
rect 583390 3304 583446 3360
<< metal3 >>
rect 293861 700770 293927 700773
rect 559649 700770 559715 700773
rect 293861 700768 559715 700770
rect 293861 700712 293866 700768
rect 293922 700712 559654 700768
rect 559710 700712 559715 700768
rect 293861 700710 559715 700712
rect 293861 700707 293927 700710
rect 559649 700707 559715 700710
rect 40493 700634 40559 700637
rect 324313 700634 324379 700637
rect 40493 700632 324379 700634
rect 40493 700576 40498 700632
rect 40554 700576 324318 700632
rect 324374 700576 324379 700632
rect 40493 700574 324379 700576
rect 40493 700571 40559 700574
rect 324313 700571 324379 700574
rect 24301 700498 24367 700501
rect 319437 700498 319503 700501
rect 24301 700496 319503 700498
rect 24301 700440 24306 700496
rect 24362 700440 319442 700496
rect 319498 700440 319503 700496
rect 24301 700438 319503 700440
rect 24301 700435 24367 700438
rect 319437 700435 319503 700438
rect 8109 700362 8175 700365
rect 325693 700362 325759 700365
rect 8109 700360 325759 700362
rect 8109 700304 8114 700360
rect 8170 700304 325698 700360
rect 325754 700304 325759 700360
rect 8109 700302 325759 700304
rect 8109 700299 8175 700302
rect 325693 700299 325759 700302
rect -960 697220 480 697460
rect 580165 697234 580231 697237
rect 583520 697234 584960 697324
rect 580165 697232 584960 697234
rect 580165 697176 580170 697232
rect 580226 697176 584960 697232
rect 580165 697174 584960 697176
rect 580165 697171 580231 697174
rect 583520 697084 584960 697174
rect -960 684314 480 684404
rect 3417 684314 3483 684317
rect -960 684312 3483 684314
rect -960 684256 3422 684312
rect 3478 684256 3483 684312
rect -960 684254 3483 684256
rect -960 684164 480 684254
rect 3417 684251 3483 684254
rect 580165 683906 580231 683909
rect 583520 683906 584960 683996
rect 580165 683904 584960 683906
rect 580165 683848 580170 683904
rect 580226 683848 584960 683904
rect 580165 683846 584960 683848
rect 580165 683843 580231 683846
rect 583520 683756 584960 683846
rect -960 671258 480 671348
rect 3509 671258 3575 671261
rect -960 671256 3575 671258
rect -960 671200 3514 671256
rect 3570 671200 3575 671256
rect -960 671198 3575 671200
rect -960 671108 480 671198
rect 3509 671195 3575 671198
rect 580165 670714 580231 670717
rect 583520 670714 584960 670804
rect 580165 670712 584960 670714
rect 580165 670656 580170 670712
rect 580226 670656 584960 670712
rect 580165 670654 584960 670656
rect 580165 670651 580231 670654
rect 583520 670564 584960 670654
rect -960 658202 480 658292
rect 3417 658202 3483 658205
rect -960 658200 3483 658202
rect -960 658144 3422 658200
rect 3478 658144 3483 658200
rect -960 658142 3483 658144
rect -960 658052 480 658142
rect 3417 658139 3483 658142
rect 583520 657236 584960 657476
rect -960 644996 480 645236
rect 580165 644058 580231 644061
rect 583520 644058 584960 644148
rect 580165 644056 584960 644058
rect 580165 644000 580170 644056
rect 580226 644000 584960 644056
rect 580165 643998 584960 644000
rect 580165 643995 580231 643998
rect 583520 643908 584960 643998
rect -960 632090 480 632180
rect 3417 632090 3483 632093
rect -960 632088 3483 632090
rect -960 632032 3422 632088
rect 3478 632032 3483 632088
rect -960 632030 3483 632032
rect -960 631940 480 632030
rect 3417 632027 3483 632030
rect 580165 630866 580231 630869
rect 583520 630866 584960 630956
rect 580165 630864 584960 630866
rect 580165 630808 580170 630864
rect 580226 630808 584960 630864
rect 580165 630806 584960 630808
rect 580165 630803 580231 630806
rect 583520 630716 584960 630806
rect -960 619170 480 619260
rect 3141 619170 3207 619173
rect -960 619168 3207 619170
rect -960 619112 3146 619168
rect 3202 619112 3207 619168
rect -960 619110 3207 619112
rect -960 619020 480 619110
rect 3141 619107 3207 619110
rect 580165 617538 580231 617541
rect 583520 617538 584960 617628
rect 580165 617536 584960 617538
rect 580165 617480 580170 617536
rect 580226 617480 584960 617536
rect 580165 617478 584960 617480
rect 580165 617475 580231 617478
rect 583520 617388 584960 617478
rect -960 606114 480 606204
rect 3233 606114 3299 606117
rect -960 606112 3299 606114
rect -960 606056 3238 606112
rect 3294 606056 3299 606112
rect -960 606054 3299 606056
rect -960 605964 480 606054
rect 3233 606051 3299 606054
rect 583520 604060 584960 604300
rect -960 592908 480 593148
rect 579797 591018 579863 591021
rect 583520 591018 584960 591108
rect 579797 591016 584960 591018
rect 579797 590960 579802 591016
rect 579858 590960 584960 591016
rect 579797 590958 584960 590960
rect 579797 590955 579863 590958
rect 583520 590868 584960 590958
rect -960 580002 480 580092
rect 3325 580002 3391 580005
rect -960 580000 3391 580002
rect -960 579944 3330 580000
rect 3386 579944 3391 580000
rect -960 579942 3391 579944
rect -960 579852 480 579942
rect 3325 579939 3391 579942
rect 580165 577690 580231 577693
rect 583520 577690 584960 577780
rect 580165 577688 584960 577690
rect 580165 577632 580170 577688
rect 580226 577632 584960 577688
rect 580165 577630 584960 577632
rect 580165 577627 580231 577630
rect 583520 577540 584960 577630
rect -960 566946 480 567036
rect 3417 566946 3483 566949
rect -960 566944 3483 566946
rect -960 566888 3422 566944
rect 3478 566888 3483 566944
rect -960 566886 3483 566888
rect -960 566796 480 566886
rect 3417 566883 3483 566886
rect 579797 564362 579863 564365
rect 583520 564362 584960 564452
rect 579797 564360 584960 564362
rect 579797 564304 579802 564360
rect 579858 564304 584960 564360
rect 579797 564302 584960 564304
rect 579797 564299 579863 564302
rect 583520 564212 584960 564302
rect -960 553890 480 553980
rect 3417 553890 3483 553893
rect -960 553888 3483 553890
rect -960 553832 3422 553888
rect 3478 553832 3483 553888
rect -960 553830 3483 553832
rect -960 553740 480 553830
rect 3417 553827 3483 553830
rect 583520 551020 584960 551260
rect -960 540684 480 540924
rect 580165 537842 580231 537845
rect 583520 537842 584960 537932
rect 580165 537840 584960 537842
rect 580165 537784 580170 537840
rect 580226 537784 584960 537840
rect 580165 537782 584960 537784
rect 580165 537779 580231 537782
rect 583520 537692 584960 537782
rect -960 527914 480 528004
rect 3417 527914 3483 527917
rect -960 527912 3483 527914
rect -960 527856 3422 527912
rect 3478 527856 3483 527912
rect -960 527854 3483 527856
rect -960 527764 480 527854
rect 3417 527851 3483 527854
rect 580165 524514 580231 524517
rect 583520 524514 584960 524604
rect 580165 524512 584960 524514
rect 580165 524456 580170 524512
rect 580226 524456 584960 524512
rect 580165 524454 584960 524456
rect 580165 524451 580231 524454
rect 583520 524364 584960 524454
rect -960 514858 480 514948
rect 3417 514858 3483 514861
rect -960 514856 3483 514858
rect -960 514800 3422 514856
rect 3478 514800 3483 514856
rect -960 514798 3483 514800
rect -960 514708 480 514798
rect 3417 514795 3483 514798
rect 580165 511322 580231 511325
rect 583520 511322 584960 511412
rect 580165 511320 584960 511322
rect 580165 511264 580170 511320
rect 580226 511264 584960 511320
rect 580165 511262 584960 511264
rect 580165 511259 580231 511262
rect 583520 511172 584960 511262
rect -960 501802 480 501892
rect 3049 501802 3115 501805
rect -960 501800 3115 501802
rect -960 501744 3054 501800
rect 3110 501744 3115 501800
rect -960 501742 3115 501744
rect -960 501652 480 501742
rect 3049 501739 3115 501742
rect 583520 497844 584960 498084
rect 242433 490242 242499 490245
rect 385677 490242 385743 490245
rect 242433 490240 385743 490242
rect 242433 490184 242438 490240
rect 242494 490184 385682 490240
rect 385738 490184 385743 490240
rect 242433 490182 385743 490184
rect 242433 490179 242499 490182
rect 385677 490179 385743 490182
rect 238569 490106 238635 490109
rect 384297 490106 384363 490109
rect 238569 490104 384363 490106
rect 238569 490048 238574 490104
rect 238630 490048 384302 490104
rect 384358 490048 384363 490104
rect 238569 490046 384363 490048
rect 238569 490043 238635 490046
rect 384297 490043 384363 490046
rect 237281 489970 237347 489973
rect 384481 489970 384547 489973
rect 237281 489968 384547 489970
rect 237281 489912 237286 489968
rect 237342 489912 384486 489968
rect 384542 489912 384547 489968
rect 237281 489910 384547 489912
rect 237281 489907 237347 489910
rect 384481 489907 384547 489910
rect -960 488596 480 488836
rect 373901 487114 373967 487117
rect 354630 487112 373967 487114
rect 354630 487056 373906 487112
rect 373962 487056 373967 487112
rect 354630 487054 373967 487056
rect 8017 486162 8083 486165
rect 354630 486162 354690 487054
rect 373901 487051 373967 487054
rect 372613 486978 372679 486981
rect 377581 486978 377647 486981
rect 8017 486160 354690 486162
rect 8017 486104 8022 486160
rect 8078 486104 354690 486160
rect 8017 486102 354690 486104
rect 368430 486976 372679 486978
rect 368430 486920 372618 486976
rect 372674 486920 372679 486976
rect 368430 486918 372679 486920
rect 8017 486099 8083 486102
rect 6177 486026 6243 486029
rect 368430 486026 368490 486918
rect 372613 486915 372679 486918
rect 373950 486976 377647 486978
rect 373950 486920 377586 486976
rect 377642 486920 377647 486976
rect 373950 486918 377647 486920
rect 6177 486024 368490 486026
rect 6177 485968 6182 486024
rect 6238 485968 368490 486024
rect 6177 485966 368490 485968
rect 6177 485963 6243 485966
rect 7833 485890 7899 485893
rect 373950 485890 374010 486918
rect 377581 486915 377647 486918
rect 7833 485888 374010 485890
rect 7833 485832 7838 485888
rect 7894 485832 374010 485888
rect 7833 485830 374010 485832
rect 7833 485827 7899 485830
rect 580165 484666 580231 484669
rect 583520 484666 584960 484756
rect 580165 484664 584960 484666
rect 580165 484608 580170 484664
rect 580226 484608 584960 484664
rect 580165 484606 584960 484608
rect 580165 484603 580231 484606
rect 583520 484516 584960 484606
rect -960 475690 480 475780
rect 2773 475690 2839 475693
rect -960 475688 2839 475690
rect -960 475632 2778 475688
rect 2834 475632 2839 475688
rect -960 475630 2839 475632
rect -960 475540 480 475630
rect 2773 475627 2839 475630
rect 580165 471474 580231 471477
rect 583520 471474 584960 471564
rect 580165 471472 584960 471474
rect 580165 471416 580170 471472
rect 580226 471416 584960 471472
rect 580165 471414 584960 471416
rect 580165 471411 580231 471414
rect 583520 471324 584960 471414
rect -960 462634 480 462724
rect 3233 462634 3299 462637
rect -960 462632 3299 462634
rect -960 462576 3238 462632
rect 3294 462576 3299 462632
rect -960 462574 3299 462576
rect -960 462484 480 462574
rect 3233 462571 3299 462574
rect 580165 458146 580231 458149
rect 583520 458146 584960 458236
rect 580165 458144 584960 458146
rect 580165 458088 580170 458144
rect 580226 458088 584960 458144
rect 580165 458086 584960 458088
rect 580165 458083 580231 458086
rect 583520 457996 584960 458086
rect -960 449578 480 449668
rect 3233 449578 3299 449581
rect -960 449576 3299 449578
rect -960 449520 3238 449576
rect 3294 449520 3299 449576
rect -960 449518 3299 449520
rect -960 449428 480 449518
rect 3233 449515 3299 449518
rect 583520 444668 584960 444908
rect -960 436508 480 436748
rect 580165 431626 580231 431629
rect 583520 431626 584960 431716
rect 580165 431624 584960 431626
rect 580165 431568 580170 431624
rect 580226 431568 584960 431624
rect 580165 431566 584960 431568
rect 580165 431563 580231 431566
rect 583520 431476 584960 431566
rect -960 423602 480 423692
rect 2773 423602 2839 423605
rect -960 423600 2839 423602
rect -960 423544 2778 423600
rect 2834 423544 2839 423600
rect -960 423542 2839 423544
rect -960 423452 480 423542
rect 2773 423539 2839 423542
rect 580165 418298 580231 418301
rect 583520 418298 584960 418388
rect 580165 418296 584960 418298
rect 580165 418240 580170 418296
rect 580226 418240 584960 418296
rect 580165 418238 584960 418240
rect 580165 418235 580231 418238
rect 583520 418148 584960 418238
rect -960 410546 480 410636
rect 3325 410546 3391 410549
rect -960 410544 3391 410546
rect -960 410488 3330 410544
rect 3386 410488 3391 410544
rect -960 410486 3391 410488
rect -960 410396 480 410486
rect 3325 410483 3391 410486
rect 580165 404970 580231 404973
rect 583520 404970 584960 405060
rect 580165 404968 584960 404970
rect 580165 404912 580170 404968
rect 580226 404912 584960 404968
rect 580165 404910 584960 404912
rect 580165 404907 580231 404910
rect 583520 404820 584960 404910
rect -960 397490 480 397580
rect 2773 397490 2839 397493
rect -960 397488 2839 397490
rect -960 397432 2778 397488
rect 2834 397432 2839 397488
rect -960 397430 2839 397432
rect -960 397340 480 397430
rect 2773 397427 2839 397430
rect 583520 391628 584960 391868
rect -960 384284 480 384524
rect 579981 378450 580047 378453
rect 583520 378450 584960 378540
rect 579981 378448 584960 378450
rect 579981 378392 579986 378448
rect 580042 378392 584960 378448
rect 579981 378390 584960 378392
rect 579981 378387 580047 378390
rect 583520 378300 584960 378390
rect -960 371378 480 371468
rect 2773 371378 2839 371381
rect -960 371376 2839 371378
rect -960 371320 2778 371376
rect 2834 371320 2839 371376
rect -960 371318 2839 371320
rect -960 371228 480 371318
rect 2773 371315 2839 371318
rect 580901 365122 580967 365125
rect 583520 365122 584960 365212
rect 580901 365120 584960 365122
rect 580901 365064 580906 365120
rect 580962 365064 584960 365120
rect 580901 365062 584960 365064
rect 580901 365059 580967 365062
rect 583520 364972 584960 365062
rect -960 358458 480 358548
rect 4061 358458 4127 358461
rect -960 358456 4127 358458
rect -960 358400 4066 358456
rect 4122 358400 4127 358456
rect -960 358398 4127 358400
rect -960 358308 480 358398
rect 4061 358395 4127 358398
rect 580165 351930 580231 351933
rect 583520 351930 584960 352020
rect 580165 351928 584960 351930
rect 580165 351872 580170 351928
rect 580226 351872 584960 351928
rect 580165 351870 584960 351872
rect 580165 351867 580231 351870
rect 583520 351780 584960 351870
rect -960 345402 480 345492
rect 3969 345402 4035 345405
rect -960 345400 4035 345402
rect -960 345344 3974 345400
rect 4030 345344 4035 345400
rect -960 345342 4035 345344
rect -960 345252 480 345342
rect 3969 345339 4035 345342
rect 583520 338452 584960 338692
rect 377857 336426 377923 336429
rect 418797 336426 418863 336429
rect 377857 336424 418863 336426
rect 377857 336368 377862 336424
rect 377918 336368 418802 336424
rect 418858 336368 418863 336424
rect 377857 336366 418863 336368
rect 377857 336363 377923 336366
rect 418797 336363 418863 336366
rect 12341 336290 12407 336293
rect 237649 336290 237715 336293
rect 12341 336288 237715 336290
rect 12341 336232 12346 336288
rect 12402 336232 237654 336288
rect 237710 336232 237715 336288
rect 12341 336230 237715 336232
rect 12341 336227 12407 336230
rect 237649 336227 237715 336230
rect 381537 336290 381603 336293
rect 422937 336290 423003 336293
rect 381537 336288 423003 336290
rect 381537 336232 381542 336288
rect 381598 336232 422942 336288
rect 422998 336232 423003 336288
rect 381537 336230 423003 336232
rect 381537 336227 381603 336230
rect 422937 336227 423003 336230
rect 10961 336154 11027 336157
rect 237373 336154 237439 336157
rect 10961 336152 237439 336154
rect 10961 336096 10966 336152
rect 11022 336096 237378 336152
rect 237434 336096 237439 336152
rect 10961 336094 237439 336096
rect 10961 336091 11027 336094
rect 237373 336091 237439 336094
rect 379697 336154 379763 336157
rect 425789 336154 425855 336157
rect 379697 336152 425855 336154
rect 379697 336096 379702 336152
rect 379758 336096 425794 336152
rect 425850 336096 425855 336152
rect 379697 336094 425855 336096
rect 379697 336091 379763 336094
rect 425789 336091 425855 336094
rect 5441 336018 5507 336021
rect 236085 336018 236151 336021
rect 5441 336016 236151 336018
rect 5441 335960 5446 336016
rect 5502 335960 236090 336016
rect 236146 335960 236151 336016
rect 5441 335958 236151 335960
rect 5441 335955 5507 335958
rect 236085 335955 236151 335958
rect 382089 336018 382155 336021
rect 451917 336018 451983 336021
rect 382089 336016 451983 336018
rect 382089 335960 382094 336016
rect 382150 335960 451922 336016
rect 451978 335960 451983 336016
rect 382089 335958 451983 335960
rect 382089 335955 382155 335958
rect 451917 335955 451983 335958
rect -960 332196 480 332436
rect 332225 330578 332291 330581
rect 332409 330578 332475 330581
rect 332225 330576 332475 330578
rect 332225 330520 332230 330576
rect 332286 330520 332414 330576
rect 332470 330520 332475 330576
rect 332225 330518 332475 330520
rect 332225 330515 332291 330518
rect 332409 330515 332475 330518
rect 580809 325274 580875 325277
rect 583520 325274 584960 325364
rect 580809 325272 584960 325274
rect 580809 325216 580814 325272
rect 580870 325216 584960 325272
rect 580809 325214 584960 325216
rect 580809 325211 580875 325214
rect 583520 325124 584960 325214
rect -960 319290 480 319380
rect 2773 319290 2839 319293
rect -960 319288 2839 319290
rect -960 319232 2778 319288
rect 2834 319232 2839 319288
rect -960 319230 2839 319232
rect -960 319140 480 319230
rect 2773 319227 2839 319230
rect 580717 312082 580783 312085
rect 583520 312082 584960 312172
rect 580717 312080 584960 312082
rect 580717 312024 580722 312080
rect 580778 312024 584960 312080
rect 580717 312022 584960 312024
rect 580717 312019 580783 312022
rect 583520 311932 584960 312022
rect -960 306234 480 306324
rect 3877 306234 3943 306237
rect -960 306232 3943 306234
rect -960 306176 3882 306232
rect 3938 306176 3943 306232
rect -960 306174 3943 306176
rect -960 306084 480 306174
rect 3877 306171 3943 306174
rect 580165 298754 580231 298757
rect 583520 298754 584960 298844
rect 580165 298752 584960 298754
rect 580165 298696 580170 298752
rect 580226 298696 584960 298752
rect 580165 298694 584960 298696
rect 580165 298691 580231 298694
rect 583520 298604 584960 298694
rect -960 293178 480 293268
rect 3141 293178 3207 293181
rect -960 293176 3207 293178
rect -960 293120 3146 293176
rect 3202 293120 3207 293176
rect -960 293118 3207 293120
rect -960 293028 480 293118
rect 3141 293115 3207 293118
rect 583520 285276 584960 285516
rect -960 279972 480 280212
rect 580165 272234 580231 272237
rect 583520 272234 584960 272324
rect 580165 272232 584960 272234
rect 580165 272176 580170 272232
rect 580226 272176 584960 272232
rect 580165 272174 584960 272176
rect 580165 272171 580231 272174
rect 583520 272084 584960 272174
rect -960 267202 480 267292
rect 2773 267202 2839 267205
rect -960 267200 2839 267202
rect -960 267144 2778 267200
rect 2834 267144 2839 267200
rect -960 267142 2839 267144
rect -960 267052 480 267142
rect 2773 267139 2839 267142
rect 580625 258906 580691 258909
rect 583520 258906 584960 258996
rect 580625 258904 584960 258906
rect 580625 258848 580630 258904
rect 580686 258848 584960 258904
rect 580625 258846 584960 258848
rect 580625 258843 580691 258846
rect 583520 258756 584960 258846
rect -960 254146 480 254236
rect 3785 254146 3851 254149
rect -960 254144 3851 254146
rect -960 254088 3790 254144
rect 3846 254088 3851 254144
rect -960 254086 3851 254088
rect -960 253996 480 254086
rect 3785 254083 3851 254086
rect 580165 245578 580231 245581
rect 583520 245578 584960 245668
rect 580165 245576 584960 245578
rect 580165 245520 580170 245576
rect 580226 245520 584960 245576
rect 580165 245518 584960 245520
rect 580165 245515 580231 245518
rect 583520 245428 584960 245518
rect -960 241090 480 241180
rect 3233 241090 3299 241093
rect -960 241088 3299 241090
rect -960 241032 3238 241088
rect 3294 241032 3299 241088
rect -960 241030 3299 241032
rect -960 240940 480 241030
rect 3233 241027 3299 241030
rect 579981 232386 580047 232389
rect 583520 232386 584960 232476
rect 579981 232384 584960 232386
rect 579981 232328 579986 232384
rect 580042 232328 584960 232384
rect 579981 232326 584960 232328
rect 579981 232323 580047 232326
rect 583520 232236 584960 232326
rect -960 227884 480 228124
rect 580533 219058 580599 219061
rect 583520 219058 584960 219148
rect 580533 219056 584960 219058
rect 580533 219000 580538 219056
rect 580594 219000 584960 219056
rect 580533 218998 584960 219000
rect 580533 218995 580599 218998
rect 583520 218908 584960 218998
rect -960 214978 480 215068
rect 3693 214978 3759 214981
rect -960 214976 3759 214978
rect -960 214920 3698 214976
rect 3754 214920 3759 214976
rect -960 214918 3759 214920
rect -960 214828 480 214918
rect 3693 214915 3759 214918
rect 580165 205730 580231 205733
rect 583520 205730 584960 205820
rect 580165 205728 584960 205730
rect 580165 205672 580170 205728
rect 580226 205672 584960 205728
rect 580165 205670 584960 205672
rect 580165 205667 580231 205670
rect 583520 205580 584960 205670
rect -960 201922 480 202012
rect 3601 201922 3667 201925
rect -960 201920 3667 201922
rect -960 201864 3606 201920
rect 3662 201864 3667 201920
rect -960 201862 3667 201864
rect -960 201772 480 201862
rect 3601 201859 3667 201862
rect 580165 192538 580231 192541
rect 583520 192538 584960 192628
rect 580165 192536 584960 192538
rect 580165 192480 580170 192536
rect 580226 192480 584960 192536
rect 580165 192478 584960 192480
rect 580165 192475 580231 192478
rect 583520 192388 584960 192478
rect -960 188866 480 188956
rect 3233 188866 3299 188869
rect -960 188864 3299 188866
rect -960 188808 3238 188864
rect 3294 188808 3299 188864
rect -960 188806 3299 188808
rect -960 188716 480 188806
rect 3233 188803 3299 188806
rect 580441 179210 580507 179213
rect 583520 179210 584960 179300
rect 580441 179208 584960 179210
rect 580441 179152 580446 179208
rect 580502 179152 584960 179208
rect 580441 179150 584960 179152
rect 580441 179147 580507 179150
rect 583520 179060 584960 179150
rect -960 175796 480 176036
rect 580165 165882 580231 165885
rect 583520 165882 584960 165972
rect 580165 165880 584960 165882
rect 580165 165824 580170 165880
rect 580226 165824 584960 165880
rect 580165 165822 584960 165824
rect 580165 165819 580231 165822
rect 583520 165732 584960 165822
rect -960 162890 480 162980
rect 3509 162890 3575 162893
rect -960 162888 3575 162890
rect -960 162832 3514 162888
rect 3570 162832 3575 162888
rect -960 162830 3575 162832
rect -960 162740 480 162830
rect 3509 162827 3575 162830
rect 579613 152690 579679 152693
rect 583520 152690 584960 152780
rect 579613 152688 584960 152690
rect 579613 152632 579618 152688
rect 579674 152632 584960 152688
rect 579613 152630 584960 152632
rect 579613 152627 579679 152630
rect 583520 152540 584960 152630
rect -960 149834 480 149924
rect 3417 149834 3483 149837
rect -960 149832 3483 149834
rect -960 149776 3422 149832
rect 3478 149776 3483 149832
rect -960 149774 3483 149776
rect -960 149684 480 149774
rect 3417 149771 3483 149774
rect 580349 139362 580415 139365
rect 583520 139362 584960 139452
rect 580349 139360 584960 139362
rect 580349 139304 580354 139360
rect 580410 139304 584960 139360
rect 580349 139302 584960 139304
rect 580349 139299 580415 139302
rect 583520 139212 584960 139302
rect -960 136778 480 136868
rect 3233 136778 3299 136781
rect -960 136776 3299 136778
rect -960 136720 3238 136776
rect 3294 136720 3299 136776
rect -960 136718 3299 136720
rect -960 136628 480 136718
rect 3233 136715 3299 136718
rect 580165 126034 580231 126037
rect 583520 126034 584960 126124
rect 580165 126032 584960 126034
rect 580165 125976 580170 126032
rect 580226 125976 584960 126032
rect 580165 125974 584960 125976
rect 580165 125971 580231 125974
rect 583520 125884 584960 125974
rect -960 123572 480 123812
rect 580165 112842 580231 112845
rect 583520 112842 584960 112932
rect 580165 112840 584960 112842
rect 580165 112784 580170 112840
rect 580226 112784 584960 112840
rect 580165 112782 584960 112784
rect 580165 112779 580231 112782
rect 583520 112692 584960 112782
rect -960 110666 480 110756
rect 2773 110666 2839 110669
rect -960 110664 2839 110666
rect -960 110608 2778 110664
rect 2834 110608 2839 110664
rect -960 110606 2839 110608
rect -960 110516 480 110606
rect 2773 110603 2839 110606
rect 580257 99514 580323 99517
rect 583520 99514 584960 99604
rect 580257 99512 584960 99514
rect 580257 99456 580262 99512
rect 580318 99456 584960 99512
rect 580257 99454 584960 99456
rect 580257 99451 580323 99454
rect 583520 99364 584960 99454
rect -960 97610 480 97700
rect 3325 97610 3391 97613
rect -960 97608 3391 97610
rect -960 97552 3330 97608
rect 3386 97552 3391 97608
rect -960 97550 3391 97552
rect -960 97460 480 97550
rect 3325 97547 3391 97550
rect 580165 86186 580231 86189
rect 583520 86186 584960 86276
rect 580165 86184 584960 86186
rect 580165 86128 580170 86184
rect 580226 86128 584960 86184
rect 580165 86126 584960 86128
rect 580165 86123 580231 86126
rect 583520 86036 584960 86126
rect -960 84690 480 84780
rect 2773 84690 2839 84693
rect -960 84688 2839 84690
rect -960 84632 2778 84688
rect 2834 84632 2839 84688
rect -960 84630 2839 84632
rect -960 84540 480 84630
rect 2773 84627 2839 84630
rect 580165 72994 580231 72997
rect 583520 72994 584960 73084
rect 580165 72992 584960 72994
rect 580165 72936 580170 72992
rect 580226 72936 584960 72992
rect 580165 72934 584960 72936
rect 580165 72931 580231 72934
rect 583520 72844 584960 72934
rect -960 71634 480 71724
rect 2773 71634 2839 71637
rect -960 71632 2839 71634
rect -960 71576 2778 71632
rect 2834 71576 2839 71632
rect -960 71574 2839 71576
rect -960 71484 480 71574
rect 2773 71571 2839 71574
rect 580165 59666 580231 59669
rect 583520 59666 584960 59756
rect 580165 59664 584960 59666
rect 580165 59608 580170 59664
rect 580226 59608 584960 59664
rect 580165 59606 584960 59608
rect 580165 59603 580231 59606
rect 583520 59516 584960 59606
rect -960 58578 480 58668
rect 3049 58578 3115 58581
rect -960 58576 3115 58578
rect -960 58520 3054 58576
rect 3110 58520 3115 58576
rect -960 58518 3115 58520
rect -960 58428 480 58518
rect 3049 58515 3115 58518
rect 580165 46338 580231 46341
rect 583520 46338 584960 46428
rect 580165 46336 584960 46338
rect 580165 46280 580170 46336
rect 580226 46280 584960 46336
rect 580165 46278 584960 46280
rect 580165 46275 580231 46278
rect 583520 46188 584960 46278
rect -960 45522 480 45612
rect 3417 45522 3483 45525
rect -960 45520 3483 45522
rect -960 45464 3422 45520
rect 3478 45464 3483 45520
rect -960 45462 3483 45464
rect -960 45372 480 45462
rect 3417 45459 3483 45462
rect 580165 33146 580231 33149
rect 583520 33146 584960 33236
rect 580165 33144 584960 33146
rect 580165 33088 580170 33144
rect 580226 33088 584960 33144
rect 580165 33086 584960 33088
rect 580165 33083 580231 33086
rect 583520 32996 584960 33086
rect -960 32466 480 32556
rect 2773 32466 2839 32469
rect -960 32464 2839 32466
rect -960 32408 2778 32464
rect 2834 32408 2839 32464
rect -960 32406 2839 32408
rect -960 32316 480 32406
rect 2773 32403 2839 32406
rect 579981 19818 580047 19821
rect 583520 19818 584960 19908
rect 579981 19816 584960 19818
rect 579981 19760 579986 19816
rect 580042 19760 584960 19816
rect 579981 19758 584960 19760
rect 579981 19755 580047 19758
rect 583520 19668 584960 19758
rect -960 19410 480 19500
rect 3049 19410 3115 19413
rect -960 19408 3115 19410
rect -960 19352 3054 19408
rect 3110 19352 3115 19408
rect -960 19350 3115 19352
rect -960 19260 480 19350
rect 3049 19347 3115 19350
rect 79685 12066 79751 12069
rect 254117 12066 254183 12069
rect 79685 12064 254183 12066
rect 79685 12008 79690 12064
rect 79746 12008 254122 12064
rect 254178 12008 254183 12064
rect 79685 12006 254183 12008
rect 79685 12003 79751 12006
rect 254117 12003 254183 12006
rect 81341 11930 81407 11933
rect 255497 11930 255563 11933
rect 81341 11928 255563 11930
rect 81341 11872 81346 11928
rect 81402 11872 255502 11928
rect 255558 11872 255563 11928
rect 81341 11870 255563 11872
rect 81341 11867 81407 11870
rect 255497 11867 255563 11870
rect 78581 11794 78647 11797
rect 254209 11794 254275 11797
rect 78581 11792 254275 11794
rect 78581 11736 78586 11792
rect 78642 11736 254214 11792
rect 254270 11736 254275 11792
rect 78581 11734 254275 11736
rect 78581 11731 78647 11734
rect 254209 11731 254275 11734
rect 1301 11658 1367 11661
rect 234613 11658 234679 11661
rect 1301 11656 234679 11658
rect 1301 11600 1306 11656
rect 1362 11600 234618 11656
rect 234674 11600 234679 11656
rect 1301 11598 234679 11600
rect 1301 11595 1367 11598
rect 234613 11595 234679 11598
rect 45461 10706 45527 10709
rect 245837 10706 245903 10709
rect 45461 10704 245903 10706
rect 45461 10648 45466 10704
rect 45522 10648 245842 10704
rect 245898 10648 245903 10704
rect 45461 10646 245903 10648
rect 45461 10643 45527 10646
rect 245837 10643 245903 10646
rect 377397 10706 377463 10709
rect 511257 10706 511323 10709
rect 377397 10704 511323 10706
rect 377397 10648 377402 10704
rect 377458 10648 511262 10704
rect 511318 10648 511323 10704
rect 377397 10646 511323 10648
rect 377397 10643 377463 10646
rect 511257 10643 511323 10646
rect 41321 10570 41387 10573
rect 244549 10570 244615 10573
rect 41321 10568 244615 10570
rect 41321 10512 41326 10568
rect 41382 10512 244554 10568
rect 244610 10512 244615 10568
rect 41321 10510 244615 10512
rect 41321 10507 41387 10510
rect 244549 10507 244615 10510
rect 360009 10570 360075 10573
rect 494697 10570 494763 10573
rect 360009 10568 494763 10570
rect 360009 10512 360014 10568
rect 360070 10512 494702 10568
rect 494758 10512 494763 10568
rect 360009 10510 494763 10512
rect 360009 10507 360075 10510
rect 494697 10507 494763 10510
rect 36997 10434 37063 10437
rect 244457 10434 244523 10437
rect 36997 10432 244523 10434
rect 36997 10376 37002 10432
rect 37058 10376 244462 10432
rect 244518 10376 244523 10432
rect 36997 10374 244523 10376
rect 36997 10371 37063 10374
rect 244457 10371 244523 10374
rect 361205 10434 361271 10437
rect 497089 10434 497155 10437
rect 361205 10432 497155 10434
rect 361205 10376 361210 10432
rect 361266 10376 497094 10432
rect 497150 10376 497155 10432
rect 361205 10374 497155 10376
rect 361205 10371 361271 10374
rect 497089 10371 497155 10374
rect 13537 10298 13603 10301
rect 237557 10298 237623 10301
rect 13537 10296 237623 10298
rect 13537 10240 13542 10296
rect 13598 10240 237562 10296
rect 237618 10240 237623 10296
rect 13537 10238 237623 10240
rect 13537 10235 13603 10238
rect 237557 10235 237623 10238
rect 362585 10298 362651 10301
rect 500585 10298 500651 10301
rect 362585 10296 500651 10298
rect 362585 10240 362590 10296
rect 362646 10240 500590 10296
rect 500646 10240 500651 10296
rect 362585 10238 500651 10240
rect 362585 10235 362651 10238
rect 500585 10235 500651 10238
rect 135253 9346 135319 9349
rect 269297 9346 269363 9349
rect 135253 9344 269363 9346
rect 135253 9288 135258 9344
rect 135314 9288 269302 9344
rect 269358 9288 269363 9344
rect 135253 9286 269363 9288
rect 135253 9283 135319 9286
rect 269297 9283 269363 9286
rect 131757 9210 131823 9213
rect 268009 9210 268075 9213
rect 131757 9208 268075 9210
rect 131757 9152 131762 9208
rect 131818 9152 268014 9208
rect 268070 9152 268075 9208
rect 131757 9150 268075 9152
rect 131757 9147 131823 9150
rect 268009 9147 268075 9150
rect 352925 9210 352991 9213
rect 467465 9210 467531 9213
rect 352925 9208 467531 9210
rect 352925 9152 352930 9208
rect 352986 9152 467470 9208
rect 467526 9152 467531 9208
rect 352925 9150 467531 9152
rect 352925 9147 352991 9150
rect 467465 9147 467531 9150
rect 30097 9074 30163 9077
rect 241789 9074 241855 9077
rect 30097 9072 241855 9074
rect 30097 9016 30102 9072
rect 30158 9016 241794 9072
rect 241850 9016 241855 9072
rect 30097 9014 241855 9016
rect 30097 9011 30163 9014
rect 241789 9011 241855 9014
rect 354397 9074 354463 9077
rect 471053 9074 471119 9077
rect 354397 9072 471119 9074
rect 354397 9016 354402 9072
rect 354458 9016 471058 9072
rect 471114 9016 471119 9072
rect 354397 9014 471119 9016
rect 354397 9011 354463 9014
rect 471053 9011 471119 9014
rect 26509 8938 26575 8941
rect 241697 8938 241763 8941
rect 26509 8936 241763 8938
rect 26509 8880 26514 8936
rect 26570 8880 241702 8936
rect 241758 8880 241763 8936
rect 26509 8878 241763 8880
rect 26509 8875 26575 8878
rect 241697 8875 241763 8878
rect 355961 8938 356027 8941
rect 478137 8938 478203 8941
rect 355961 8936 478203 8938
rect 355961 8880 355966 8936
rect 356022 8880 478142 8936
rect 478198 8880 478203 8936
rect 355961 8878 478203 8880
rect 355961 8875 356027 8878
rect 478137 8875 478203 8878
rect 21817 7986 21883 7989
rect 240409 7986 240475 7989
rect 21817 7984 240475 7986
rect 21817 7928 21822 7984
rect 21878 7928 240414 7984
rect 240470 7928 240475 7984
rect 21817 7926 240475 7928
rect 21817 7923 21883 7926
rect 240409 7923 240475 7926
rect 376569 7986 376635 7989
rect 559741 7986 559807 7989
rect 376569 7984 559807 7986
rect 376569 7928 376574 7984
rect 376630 7928 559746 7984
rect 559802 7928 559807 7984
rect 376569 7926 559807 7928
rect 376569 7923 376635 7926
rect 559741 7923 559807 7926
rect 17033 7850 17099 7853
rect 238937 7850 239003 7853
rect 17033 7848 239003 7850
rect 17033 7792 17038 7848
rect 17094 7792 238942 7848
rect 238998 7792 239003 7848
rect 17033 7790 239003 7792
rect 17033 7787 17099 7790
rect 238937 7787 239003 7790
rect 377857 7850 377923 7853
rect 563237 7850 563303 7853
rect 377857 7848 563303 7850
rect 377857 7792 377862 7848
rect 377918 7792 563242 7848
rect 563298 7792 563303 7848
rect 377857 7790 563303 7792
rect 377857 7787 377923 7790
rect 563237 7787 563303 7790
rect 12249 7714 12315 7717
rect 237465 7714 237531 7717
rect 12249 7712 237531 7714
rect 12249 7656 12254 7712
rect 12310 7656 237470 7712
rect 237526 7656 237531 7712
rect 12249 7654 237531 7656
rect 12249 7651 12315 7654
rect 237465 7651 237531 7654
rect 379145 7714 379211 7717
rect 570321 7714 570387 7717
rect 379145 7712 570387 7714
rect 379145 7656 379150 7712
rect 379206 7656 570326 7712
rect 570382 7656 570387 7712
rect 379145 7654 570387 7656
rect 379145 7651 379211 7654
rect 570321 7651 570387 7654
rect 8753 7578 8819 7581
rect 236177 7578 236243 7581
rect 8753 7576 236243 7578
rect 8753 7520 8758 7576
rect 8814 7520 236182 7576
rect 236238 7520 236243 7576
rect 8753 7518 236243 7520
rect 8753 7515 8819 7518
rect 236177 7515 236243 7518
rect 380617 7578 380683 7581
rect 573909 7578 573975 7581
rect 380617 7576 573975 7578
rect 380617 7520 380622 7576
rect 380678 7520 573914 7576
rect 573970 7520 573975 7576
rect 380617 7518 573975 7520
rect 380617 7515 380683 7518
rect 573909 7515 573975 7518
rect 58433 6626 58499 6629
rect 248505 6626 248571 6629
rect 58433 6624 248571 6626
rect -960 6490 480 6580
rect 58433 6568 58438 6624
rect 58494 6568 248510 6624
rect 248566 6568 248571 6624
rect 58433 6566 248571 6568
rect 58433 6563 58499 6566
rect 248505 6563 248571 6566
rect 353017 6626 353083 6629
rect 466269 6626 466335 6629
rect 353017 6624 466335 6626
rect 353017 6568 353022 6624
rect 353078 6568 466274 6624
rect 466330 6568 466335 6624
rect 353017 6566 466335 6568
rect 353017 6563 353083 6566
rect 466269 6563 466335 6566
rect 580165 6626 580231 6629
rect 583520 6626 584960 6716
rect 580165 6624 584960 6626
rect 580165 6568 580170 6624
rect 580226 6568 584960 6624
rect 580165 6566 584960 6568
rect 580165 6563 580231 6566
rect 3417 6490 3483 6493
rect -960 6488 3483 6490
rect -960 6432 3422 6488
rect 3478 6432 3483 6488
rect -960 6430 3483 6432
rect -960 6340 480 6430
rect 3417 6427 3483 6430
rect 54937 6490 55003 6493
rect 248597 6490 248663 6493
rect 54937 6488 248663 6490
rect 54937 6432 54942 6488
rect 54998 6432 248602 6488
rect 248658 6432 248663 6488
rect 54937 6430 248663 6432
rect 54937 6427 55003 6430
rect 248597 6427 248663 6430
rect 354489 6490 354555 6493
rect 469857 6490 469923 6493
rect 354489 6488 469923 6490
rect 354489 6432 354494 6488
rect 354550 6432 469862 6488
rect 469918 6432 469923 6488
rect 583520 6476 584960 6566
rect 354489 6430 469923 6432
rect 354489 6427 354555 6430
rect 469857 6427 469923 6430
rect 51349 6354 51415 6357
rect 247217 6354 247283 6357
rect 51349 6352 247283 6354
rect 51349 6296 51354 6352
rect 51410 6296 247222 6352
rect 247278 6296 247283 6352
rect 51349 6294 247283 6296
rect 51349 6291 51415 6294
rect 247217 6291 247283 6294
rect 379237 6354 379303 6357
rect 566825 6354 566891 6357
rect 379237 6352 566891 6354
rect 379237 6296 379242 6352
rect 379298 6296 566830 6352
rect 566886 6296 566891 6352
rect 379237 6294 566891 6296
rect 379237 6291 379303 6294
rect 566825 6291 566891 6294
rect 47853 6218 47919 6221
rect 247125 6218 247191 6221
rect 47853 6216 247191 6218
rect 47853 6160 47858 6216
rect 47914 6160 247130 6216
rect 247186 6160 247191 6216
rect 47853 6158 247191 6160
rect 47853 6155 47919 6158
rect 247125 6155 247191 6158
rect 382089 6218 382155 6221
rect 577405 6218 577471 6221
rect 382089 6216 577471 6218
rect 382089 6160 382094 6216
rect 382150 6160 577410 6216
rect 577466 6160 577471 6216
rect 382089 6158 577471 6160
rect 382089 6155 382155 6158
rect 577405 6155 577471 6158
rect 168373 5266 168439 5269
rect 243537 5266 243603 5269
rect 168373 5264 243603 5266
rect 168373 5208 168378 5264
rect 168434 5208 243542 5264
rect 243598 5208 243603 5264
rect 168373 5206 243603 5208
rect 168373 5203 168439 5206
rect 243537 5203 243603 5206
rect 376661 5266 376727 5269
rect 558545 5266 558611 5269
rect 376661 5264 558611 5266
rect 376661 5208 376666 5264
rect 376722 5208 558550 5264
rect 558606 5208 558611 5264
rect 376661 5206 558611 5208
rect 376661 5203 376727 5206
rect 558545 5203 558611 5206
rect 175457 5130 175523 5133
rect 278773 5130 278839 5133
rect 175457 5128 278839 5130
rect 175457 5072 175462 5128
rect 175518 5072 278778 5128
rect 278834 5072 278839 5128
rect 175457 5070 278839 5072
rect 175457 5067 175523 5070
rect 278773 5067 278839 5070
rect 377949 5130 378015 5133
rect 565629 5130 565695 5133
rect 377949 5128 565695 5130
rect 377949 5072 377954 5128
rect 378010 5072 565634 5128
rect 565690 5072 565695 5128
rect 377949 5070 565695 5072
rect 377949 5067 378015 5070
rect 565629 5067 565695 5070
rect 132953 4994 133019 4997
rect 267733 4994 267799 4997
rect 132953 4992 267799 4994
rect 132953 4936 132958 4992
rect 133014 4936 267738 4992
rect 267794 4936 267799 4992
rect 132953 4934 267799 4936
rect 132953 4931 133019 4934
rect 267733 4931 267799 4934
rect 380801 4994 380867 4997
rect 572713 4994 572779 4997
rect 380801 4992 572779 4994
rect 380801 4936 380806 4992
rect 380862 4936 572718 4992
rect 572774 4936 572779 4992
rect 380801 4934 572779 4936
rect 380801 4931 380867 4934
rect 572713 4931 572779 4934
rect 129365 4858 129431 4861
rect 266721 4858 266787 4861
rect 129365 4856 266787 4858
rect 129365 4800 129370 4856
rect 129426 4800 266726 4856
rect 266782 4800 266787 4856
rect 129365 4798 266787 4800
rect 129365 4795 129431 4798
rect 266721 4795 266787 4798
rect 380709 4858 380775 4861
rect 576301 4858 576367 4861
rect 380709 4856 576367 4858
rect 380709 4800 380714 4856
rect 380770 4800 576306 4856
rect 576362 4800 576367 4856
rect 380709 4798 576367 4800
rect 380709 4795 380775 4798
rect 576301 4795 576367 4798
rect 335261 4042 335327 4045
rect 394233 4042 394299 4045
rect 335261 4040 394299 4042
rect 335261 3984 335266 4040
rect 335322 3984 394238 4040
rect 394294 3984 394299 4040
rect 335261 3982 394299 3984
rect 335261 3979 335327 3982
rect 394233 3979 394299 3982
rect 336549 3906 336615 3909
rect 397729 3906 397795 3909
rect 336549 3904 397795 3906
rect 336549 3848 336554 3904
rect 336610 3848 397734 3904
rect 397790 3848 397795 3904
rect 336549 3846 397795 3848
rect 336549 3843 336615 3846
rect 397729 3843 397795 3846
rect 19425 3770 19491 3773
rect 238845 3770 238911 3773
rect 19425 3768 238911 3770
rect 19425 3712 19430 3768
rect 19486 3712 238850 3768
rect 238906 3712 238911 3768
rect 19425 3710 238911 3712
rect 19425 3707 19491 3710
rect 238845 3707 238911 3710
rect 267733 3770 267799 3773
rect 302509 3770 302575 3773
rect 267733 3768 302575 3770
rect 267733 3712 267738 3768
rect 267794 3712 302514 3768
rect 302570 3712 302575 3768
rect 267733 3710 302575 3712
rect 267733 3707 267799 3710
rect 302509 3707 302575 3710
rect 336641 3770 336707 3773
rect 401317 3770 401383 3773
rect 336641 3768 401383 3770
rect 336641 3712 336646 3768
rect 336702 3712 401322 3768
rect 401378 3712 401383 3768
rect 336641 3710 401383 3712
rect 336641 3707 336707 3710
rect 401317 3707 401383 3710
rect 451917 3770 451983 3773
rect 582189 3770 582255 3773
rect 451917 3768 582255 3770
rect 451917 3712 451922 3768
rect 451978 3712 582194 3768
rect 582250 3712 582255 3768
rect 451917 3710 582255 3712
rect 451917 3707 451983 3710
rect 582189 3707 582255 3710
rect 14733 3634 14799 3637
rect 237373 3634 237439 3637
rect 14733 3632 237439 3634
rect 14733 3576 14738 3632
rect 14794 3576 237378 3632
rect 237434 3576 237439 3632
rect 14733 3574 237439 3576
rect 14733 3571 14799 3574
rect 237373 3571 237439 3574
rect 260649 3634 260715 3637
rect 300945 3634 301011 3637
rect 260649 3632 301011 3634
rect 260649 3576 260654 3632
rect 260710 3576 300950 3632
rect 301006 3576 301011 3632
rect 260649 3574 301011 3576
rect 260649 3571 260715 3574
rect 300945 3571 301011 3574
rect 339401 3634 339467 3637
rect 411897 3634 411963 3637
rect 339401 3632 411963 3634
rect 339401 3576 339406 3632
rect 339462 3576 411902 3632
rect 411958 3576 411963 3632
rect 339401 3574 411963 3576
rect 339401 3571 339467 3574
rect 411897 3571 411963 3574
rect 422937 3634 423003 3637
rect 578601 3634 578667 3637
rect 422937 3632 578667 3634
rect 422937 3576 422942 3632
rect 422998 3576 578606 3632
rect 578662 3576 578667 3632
rect 422937 3574 578667 3576
rect 422937 3571 423003 3574
rect 578601 3571 578667 3574
rect 15929 3498 15995 3501
rect 239029 3498 239095 3501
rect 15929 3496 239095 3498
rect 15929 3440 15934 3496
rect 15990 3440 239034 3496
rect 239090 3440 239095 3496
rect 15929 3438 239095 3440
rect 15929 3435 15995 3438
rect 239029 3435 239095 3438
rect 240501 3498 240567 3501
rect 295425 3498 295491 3501
rect 240501 3496 295491 3498
rect 240501 3440 240506 3496
rect 240562 3440 295430 3496
rect 295486 3440 295491 3496
rect 240501 3438 295491 3440
rect 240501 3435 240567 3438
rect 295425 3435 295491 3438
rect 379421 3498 379487 3501
rect 568021 3498 568087 3501
rect 379421 3496 568087 3498
rect 379421 3440 379426 3496
rect 379482 3440 568026 3496
rect 568082 3440 568087 3496
rect 379421 3438 568087 3440
rect 379421 3435 379487 3438
rect 568021 3435 568087 3438
rect 6453 3362 6519 3365
rect 236269 3362 236335 3365
rect 6453 3360 236335 3362
rect 6453 3304 6458 3360
rect 6514 3304 236274 3360
rect 236330 3304 236335 3360
rect 6453 3302 236335 3304
rect 6453 3299 6519 3302
rect 236269 3299 236335 3302
rect 239305 3362 239371 3365
rect 295517 3362 295583 3365
rect 239305 3360 295583 3362
rect 239305 3304 239310 3360
rect 239366 3304 295522 3360
rect 295578 3304 295583 3360
rect 239305 3302 295583 3304
rect 239305 3299 239371 3302
rect 295517 3299 295583 3302
rect 382181 3362 382247 3365
rect 583385 3362 583451 3365
rect 382181 3360 583451 3362
rect 382181 3304 382186 3360
rect 382242 3304 583390 3360
rect 583446 3304 583451 3360
rect 382181 3302 583451 3304
rect 382181 3299 382247 3302
rect 583385 3299 583451 3302
<< metal4 >>
rect -8726 711558 -8106 711590
rect -8726 711002 -8694 711558
rect -8138 711002 -8106 711558
rect -8726 680614 -8106 711002
rect -8726 680058 -8694 680614
rect -8138 680058 -8106 680614
rect -8726 644614 -8106 680058
rect -8726 644058 -8694 644614
rect -8138 644058 -8106 644614
rect -8726 608614 -8106 644058
rect -8726 608058 -8694 608614
rect -8138 608058 -8106 608614
rect -8726 572614 -8106 608058
rect -8726 572058 -8694 572614
rect -8138 572058 -8106 572614
rect -8726 536614 -8106 572058
rect -8726 536058 -8694 536614
rect -8138 536058 -8106 536614
rect -8726 500614 -8106 536058
rect -8726 500058 -8694 500614
rect -8138 500058 -8106 500614
rect -8726 464614 -8106 500058
rect -8726 464058 -8694 464614
rect -8138 464058 -8106 464614
rect -8726 428614 -8106 464058
rect -8726 428058 -8694 428614
rect -8138 428058 -8106 428614
rect -8726 392614 -8106 428058
rect -8726 392058 -8694 392614
rect -8138 392058 -8106 392614
rect -8726 356614 -8106 392058
rect -8726 356058 -8694 356614
rect -8138 356058 -8106 356614
rect -8726 320614 -8106 356058
rect -8726 320058 -8694 320614
rect -8138 320058 -8106 320614
rect -8726 284614 -8106 320058
rect -8726 284058 -8694 284614
rect -8138 284058 -8106 284614
rect -8726 248614 -8106 284058
rect -8726 248058 -8694 248614
rect -8138 248058 -8106 248614
rect -8726 212614 -8106 248058
rect -8726 212058 -8694 212614
rect -8138 212058 -8106 212614
rect -8726 176614 -8106 212058
rect -8726 176058 -8694 176614
rect -8138 176058 -8106 176614
rect -8726 140614 -8106 176058
rect -8726 140058 -8694 140614
rect -8138 140058 -8106 140614
rect -8726 104614 -8106 140058
rect -8726 104058 -8694 104614
rect -8138 104058 -8106 104614
rect -8726 68614 -8106 104058
rect -8726 68058 -8694 68614
rect -8138 68058 -8106 68614
rect -8726 32614 -8106 68058
rect -8726 32058 -8694 32614
rect -8138 32058 -8106 32614
rect -8726 -7066 -8106 32058
rect -7766 710598 -7146 710630
rect -7766 710042 -7734 710598
rect -7178 710042 -7146 710598
rect -7766 698614 -7146 710042
rect 12954 710598 13574 711590
rect 12954 710042 12986 710598
rect 13542 710042 13574 710598
rect -7766 698058 -7734 698614
rect -7178 698058 -7146 698614
rect -7766 662614 -7146 698058
rect -7766 662058 -7734 662614
rect -7178 662058 -7146 662614
rect -7766 626614 -7146 662058
rect -7766 626058 -7734 626614
rect -7178 626058 -7146 626614
rect -7766 590614 -7146 626058
rect -7766 590058 -7734 590614
rect -7178 590058 -7146 590614
rect -7766 554614 -7146 590058
rect -7766 554058 -7734 554614
rect -7178 554058 -7146 554614
rect -7766 518614 -7146 554058
rect -7766 518058 -7734 518614
rect -7178 518058 -7146 518614
rect -7766 482614 -7146 518058
rect -7766 482058 -7734 482614
rect -7178 482058 -7146 482614
rect -7766 446614 -7146 482058
rect -7766 446058 -7734 446614
rect -7178 446058 -7146 446614
rect -7766 410614 -7146 446058
rect -7766 410058 -7734 410614
rect -7178 410058 -7146 410614
rect -7766 374614 -7146 410058
rect -7766 374058 -7734 374614
rect -7178 374058 -7146 374614
rect -7766 338614 -7146 374058
rect -7766 338058 -7734 338614
rect -7178 338058 -7146 338614
rect -7766 302614 -7146 338058
rect -7766 302058 -7734 302614
rect -7178 302058 -7146 302614
rect -7766 266614 -7146 302058
rect -7766 266058 -7734 266614
rect -7178 266058 -7146 266614
rect -7766 230614 -7146 266058
rect -7766 230058 -7734 230614
rect -7178 230058 -7146 230614
rect -7766 194614 -7146 230058
rect -7766 194058 -7734 194614
rect -7178 194058 -7146 194614
rect -7766 158614 -7146 194058
rect -7766 158058 -7734 158614
rect -7178 158058 -7146 158614
rect -7766 122614 -7146 158058
rect -7766 122058 -7734 122614
rect -7178 122058 -7146 122614
rect -7766 86614 -7146 122058
rect -7766 86058 -7734 86614
rect -7178 86058 -7146 86614
rect -7766 50614 -7146 86058
rect -7766 50058 -7734 50614
rect -7178 50058 -7146 50614
rect -7766 14614 -7146 50058
rect -7766 14058 -7734 14614
rect -7178 14058 -7146 14614
rect -7766 -6106 -7146 14058
rect -6806 709638 -6186 709670
rect -6806 709082 -6774 709638
rect -6218 709082 -6186 709638
rect -6806 676894 -6186 709082
rect -6806 676338 -6774 676894
rect -6218 676338 -6186 676894
rect -6806 640894 -6186 676338
rect -6806 640338 -6774 640894
rect -6218 640338 -6186 640894
rect -6806 604894 -6186 640338
rect -6806 604338 -6774 604894
rect -6218 604338 -6186 604894
rect -6806 568894 -6186 604338
rect -6806 568338 -6774 568894
rect -6218 568338 -6186 568894
rect -6806 532894 -6186 568338
rect -6806 532338 -6774 532894
rect -6218 532338 -6186 532894
rect -6806 496894 -6186 532338
rect -6806 496338 -6774 496894
rect -6218 496338 -6186 496894
rect -6806 460894 -6186 496338
rect -6806 460338 -6774 460894
rect -6218 460338 -6186 460894
rect -6806 424894 -6186 460338
rect -6806 424338 -6774 424894
rect -6218 424338 -6186 424894
rect -6806 388894 -6186 424338
rect -6806 388338 -6774 388894
rect -6218 388338 -6186 388894
rect -6806 352894 -6186 388338
rect -6806 352338 -6774 352894
rect -6218 352338 -6186 352894
rect -6806 316894 -6186 352338
rect -6806 316338 -6774 316894
rect -6218 316338 -6186 316894
rect -6806 280894 -6186 316338
rect -6806 280338 -6774 280894
rect -6218 280338 -6186 280894
rect -6806 244894 -6186 280338
rect -6806 244338 -6774 244894
rect -6218 244338 -6186 244894
rect -6806 208894 -6186 244338
rect -6806 208338 -6774 208894
rect -6218 208338 -6186 208894
rect -6806 172894 -6186 208338
rect -6806 172338 -6774 172894
rect -6218 172338 -6186 172894
rect -6806 136894 -6186 172338
rect -6806 136338 -6774 136894
rect -6218 136338 -6186 136894
rect -6806 100894 -6186 136338
rect -6806 100338 -6774 100894
rect -6218 100338 -6186 100894
rect -6806 64894 -6186 100338
rect -6806 64338 -6774 64894
rect -6218 64338 -6186 64894
rect -6806 28894 -6186 64338
rect -6806 28338 -6774 28894
rect -6218 28338 -6186 28894
rect -6806 -5146 -6186 28338
rect -5846 708678 -5226 708710
rect -5846 708122 -5814 708678
rect -5258 708122 -5226 708678
rect -5846 694894 -5226 708122
rect 9234 708678 9854 709670
rect 9234 708122 9266 708678
rect 9822 708122 9854 708678
rect -5846 694338 -5814 694894
rect -5258 694338 -5226 694894
rect -5846 658894 -5226 694338
rect -5846 658338 -5814 658894
rect -5258 658338 -5226 658894
rect -5846 622894 -5226 658338
rect -5846 622338 -5814 622894
rect -5258 622338 -5226 622894
rect -5846 586894 -5226 622338
rect -5846 586338 -5814 586894
rect -5258 586338 -5226 586894
rect -5846 550894 -5226 586338
rect -5846 550338 -5814 550894
rect -5258 550338 -5226 550894
rect -5846 514894 -5226 550338
rect -5846 514338 -5814 514894
rect -5258 514338 -5226 514894
rect -5846 478894 -5226 514338
rect -5846 478338 -5814 478894
rect -5258 478338 -5226 478894
rect -5846 442894 -5226 478338
rect -5846 442338 -5814 442894
rect -5258 442338 -5226 442894
rect -5846 406894 -5226 442338
rect -5846 406338 -5814 406894
rect -5258 406338 -5226 406894
rect -5846 370894 -5226 406338
rect -5846 370338 -5814 370894
rect -5258 370338 -5226 370894
rect -5846 334894 -5226 370338
rect -5846 334338 -5814 334894
rect -5258 334338 -5226 334894
rect -5846 298894 -5226 334338
rect -5846 298338 -5814 298894
rect -5258 298338 -5226 298894
rect -5846 262894 -5226 298338
rect -5846 262338 -5814 262894
rect -5258 262338 -5226 262894
rect -5846 226894 -5226 262338
rect -5846 226338 -5814 226894
rect -5258 226338 -5226 226894
rect -5846 190894 -5226 226338
rect -5846 190338 -5814 190894
rect -5258 190338 -5226 190894
rect -5846 154894 -5226 190338
rect -5846 154338 -5814 154894
rect -5258 154338 -5226 154894
rect -5846 118894 -5226 154338
rect -5846 118338 -5814 118894
rect -5258 118338 -5226 118894
rect -5846 82894 -5226 118338
rect -5846 82338 -5814 82894
rect -5258 82338 -5226 82894
rect -5846 46894 -5226 82338
rect -5846 46338 -5814 46894
rect -5258 46338 -5226 46894
rect -5846 10894 -5226 46338
rect -5846 10338 -5814 10894
rect -5258 10338 -5226 10894
rect -5846 -4186 -5226 10338
rect -4886 707718 -4266 707750
rect -4886 707162 -4854 707718
rect -4298 707162 -4266 707718
rect -4886 673174 -4266 707162
rect -4886 672618 -4854 673174
rect -4298 672618 -4266 673174
rect -4886 637174 -4266 672618
rect -4886 636618 -4854 637174
rect -4298 636618 -4266 637174
rect -4886 601174 -4266 636618
rect -4886 600618 -4854 601174
rect -4298 600618 -4266 601174
rect -4886 565174 -4266 600618
rect -4886 564618 -4854 565174
rect -4298 564618 -4266 565174
rect -4886 529174 -4266 564618
rect -4886 528618 -4854 529174
rect -4298 528618 -4266 529174
rect -4886 493174 -4266 528618
rect -4886 492618 -4854 493174
rect -4298 492618 -4266 493174
rect -4886 457174 -4266 492618
rect -4886 456618 -4854 457174
rect -4298 456618 -4266 457174
rect -4886 421174 -4266 456618
rect -4886 420618 -4854 421174
rect -4298 420618 -4266 421174
rect -4886 385174 -4266 420618
rect -4886 384618 -4854 385174
rect -4298 384618 -4266 385174
rect -4886 349174 -4266 384618
rect -4886 348618 -4854 349174
rect -4298 348618 -4266 349174
rect -4886 313174 -4266 348618
rect -4886 312618 -4854 313174
rect -4298 312618 -4266 313174
rect -4886 277174 -4266 312618
rect -4886 276618 -4854 277174
rect -4298 276618 -4266 277174
rect -4886 241174 -4266 276618
rect -4886 240618 -4854 241174
rect -4298 240618 -4266 241174
rect -4886 205174 -4266 240618
rect -4886 204618 -4854 205174
rect -4298 204618 -4266 205174
rect -4886 169174 -4266 204618
rect -4886 168618 -4854 169174
rect -4298 168618 -4266 169174
rect -4886 133174 -4266 168618
rect -4886 132618 -4854 133174
rect -4298 132618 -4266 133174
rect -4886 97174 -4266 132618
rect -4886 96618 -4854 97174
rect -4298 96618 -4266 97174
rect -4886 61174 -4266 96618
rect -4886 60618 -4854 61174
rect -4298 60618 -4266 61174
rect -4886 25174 -4266 60618
rect -4886 24618 -4854 25174
rect -4298 24618 -4266 25174
rect -4886 -3226 -4266 24618
rect -3926 706758 -3306 706790
rect -3926 706202 -3894 706758
rect -3338 706202 -3306 706758
rect -3926 691174 -3306 706202
rect 5514 706758 6134 707750
rect 5514 706202 5546 706758
rect 6102 706202 6134 706758
rect -3926 690618 -3894 691174
rect -3338 690618 -3306 691174
rect -3926 655174 -3306 690618
rect -3926 654618 -3894 655174
rect -3338 654618 -3306 655174
rect -3926 619174 -3306 654618
rect -3926 618618 -3894 619174
rect -3338 618618 -3306 619174
rect -3926 583174 -3306 618618
rect -3926 582618 -3894 583174
rect -3338 582618 -3306 583174
rect -3926 547174 -3306 582618
rect -3926 546618 -3894 547174
rect -3338 546618 -3306 547174
rect -3926 511174 -3306 546618
rect -3926 510618 -3894 511174
rect -3338 510618 -3306 511174
rect -3926 475174 -3306 510618
rect -3926 474618 -3894 475174
rect -3338 474618 -3306 475174
rect -3926 439174 -3306 474618
rect -3926 438618 -3894 439174
rect -3338 438618 -3306 439174
rect -3926 403174 -3306 438618
rect -3926 402618 -3894 403174
rect -3338 402618 -3306 403174
rect -3926 367174 -3306 402618
rect -3926 366618 -3894 367174
rect -3338 366618 -3306 367174
rect -3926 331174 -3306 366618
rect -3926 330618 -3894 331174
rect -3338 330618 -3306 331174
rect -3926 295174 -3306 330618
rect -3926 294618 -3894 295174
rect -3338 294618 -3306 295174
rect -3926 259174 -3306 294618
rect -3926 258618 -3894 259174
rect -3338 258618 -3306 259174
rect -3926 223174 -3306 258618
rect -3926 222618 -3894 223174
rect -3338 222618 -3306 223174
rect -3926 187174 -3306 222618
rect -3926 186618 -3894 187174
rect -3338 186618 -3306 187174
rect -3926 151174 -3306 186618
rect -3926 150618 -3894 151174
rect -3338 150618 -3306 151174
rect -3926 115174 -3306 150618
rect -3926 114618 -3894 115174
rect -3338 114618 -3306 115174
rect -3926 79174 -3306 114618
rect -3926 78618 -3894 79174
rect -3338 78618 -3306 79174
rect -3926 43174 -3306 78618
rect -3926 42618 -3894 43174
rect -3338 42618 -3306 43174
rect -3926 7174 -3306 42618
rect -3926 6618 -3894 7174
rect -3338 6618 -3306 7174
rect -3926 -2266 -3306 6618
rect -2966 705798 -2346 705830
rect -2966 705242 -2934 705798
rect -2378 705242 -2346 705798
rect -2966 669454 -2346 705242
rect -2966 668898 -2934 669454
rect -2378 668898 -2346 669454
rect -2966 633454 -2346 668898
rect -2966 632898 -2934 633454
rect -2378 632898 -2346 633454
rect -2966 597454 -2346 632898
rect -2966 596898 -2934 597454
rect -2378 596898 -2346 597454
rect -2966 561454 -2346 596898
rect -2966 560898 -2934 561454
rect -2378 560898 -2346 561454
rect -2966 525454 -2346 560898
rect -2966 524898 -2934 525454
rect -2378 524898 -2346 525454
rect -2966 489454 -2346 524898
rect -2966 488898 -2934 489454
rect -2378 488898 -2346 489454
rect -2966 453454 -2346 488898
rect -2966 452898 -2934 453454
rect -2378 452898 -2346 453454
rect -2966 417454 -2346 452898
rect -2966 416898 -2934 417454
rect -2378 416898 -2346 417454
rect -2966 381454 -2346 416898
rect -2966 380898 -2934 381454
rect -2378 380898 -2346 381454
rect -2966 345454 -2346 380898
rect -2966 344898 -2934 345454
rect -2378 344898 -2346 345454
rect -2966 309454 -2346 344898
rect -2966 308898 -2934 309454
rect -2378 308898 -2346 309454
rect -2966 273454 -2346 308898
rect -2966 272898 -2934 273454
rect -2378 272898 -2346 273454
rect -2966 237454 -2346 272898
rect -2966 236898 -2934 237454
rect -2378 236898 -2346 237454
rect -2966 201454 -2346 236898
rect -2966 200898 -2934 201454
rect -2378 200898 -2346 201454
rect -2966 165454 -2346 200898
rect -2966 164898 -2934 165454
rect -2378 164898 -2346 165454
rect -2966 129454 -2346 164898
rect -2966 128898 -2934 129454
rect -2378 128898 -2346 129454
rect -2966 93454 -2346 128898
rect -2966 92898 -2934 93454
rect -2378 92898 -2346 93454
rect -2966 57454 -2346 92898
rect -2966 56898 -2934 57454
rect -2378 56898 -2346 57454
rect -2966 21454 -2346 56898
rect -2966 20898 -2934 21454
rect -2378 20898 -2346 21454
rect -2966 -1306 -2346 20898
rect -2006 704838 -1386 704870
rect -2006 704282 -1974 704838
rect -1418 704282 -1386 704838
rect -2006 687454 -1386 704282
rect -2006 686898 -1974 687454
rect -1418 686898 -1386 687454
rect -2006 651454 -1386 686898
rect -2006 650898 -1974 651454
rect -1418 650898 -1386 651454
rect -2006 615454 -1386 650898
rect -2006 614898 -1974 615454
rect -1418 614898 -1386 615454
rect -2006 579454 -1386 614898
rect -2006 578898 -1974 579454
rect -1418 578898 -1386 579454
rect -2006 543454 -1386 578898
rect -2006 542898 -1974 543454
rect -1418 542898 -1386 543454
rect -2006 507454 -1386 542898
rect -2006 506898 -1974 507454
rect -1418 506898 -1386 507454
rect -2006 471454 -1386 506898
rect -2006 470898 -1974 471454
rect -1418 470898 -1386 471454
rect -2006 435454 -1386 470898
rect -2006 434898 -1974 435454
rect -1418 434898 -1386 435454
rect -2006 399454 -1386 434898
rect -2006 398898 -1974 399454
rect -1418 398898 -1386 399454
rect -2006 363454 -1386 398898
rect -2006 362898 -1974 363454
rect -1418 362898 -1386 363454
rect -2006 327454 -1386 362898
rect -2006 326898 -1974 327454
rect -1418 326898 -1386 327454
rect -2006 291454 -1386 326898
rect -2006 290898 -1974 291454
rect -1418 290898 -1386 291454
rect -2006 255454 -1386 290898
rect -2006 254898 -1974 255454
rect -1418 254898 -1386 255454
rect -2006 219454 -1386 254898
rect -2006 218898 -1974 219454
rect -1418 218898 -1386 219454
rect -2006 183454 -1386 218898
rect -2006 182898 -1974 183454
rect -1418 182898 -1386 183454
rect -2006 147454 -1386 182898
rect -2006 146898 -1974 147454
rect -1418 146898 -1386 147454
rect -2006 111454 -1386 146898
rect -2006 110898 -1974 111454
rect -1418 110898 -1386 111454
rect -2006 75454 -1386 110898
rect -2006 74898 -1974 75454
rect -1418 74898 -1386 75454
rect -2006 39454 -1386 74898
rect -2006 38898 -1974 39454
rect -1418 38898 -1386 39454
rect -2006 3454 -1386 38898
rect -2006 2898 -1974 3454
rect -1418 2898 -1386 3454
rect -2006 -346 -1386 2898
rect -2006 -902 -1974 -346
rect -1418 -902 -1386 -346
rect -2006 -934 -1386 -902
rect 1794 704838 2414 705830
rect 1794 704282 1826 704838
rect 2382 704282 2414 704838
rect 1794 687454 2414 704282
rect 1794 686898 1826 687454
rect 2382 686898 2414 687454
rect 1794 651454 2414 686898
rect 1794 650898 1826 651454
rect 2382 650898 2414 651454
rect 1794 615454 2414 650898
rect 1794 614898 1826 615454
rect 2382 614898 2414 615454
rect 1794 579454 2414 614898
rect 1794 578898 1826 579454
rect 2382 578898 2414 579454
rect 1794 543454 2414 578898
rect 1794 542898 1826 543454
rect 2382 542898 2414 543454
rect 1794 507454 2414 542898
rect 1794 506898 1826 507454
rect 2382 506898 2414 507454
rect 1794 471454 2414 506898
rect 1794 470898 1826 471454
rect 2382 470898 2414 471454
rect 1794 435454 2414 470898
rect 1794 434898 1826 435454
rect 2382 434898 2414 435454
rect 1794 399454 2414 434898
rect 1794 398898 1826 399454
rect 2382 398898 2414 399454
rect 1794 363454 2414 398898
rect 1794 362898 1826 363454
rect 2382 362898 2414 363454
rect 1794 327454 2414 362898
rect 1794 326898 1826 327454
rect 2382 326898 2414 327454
rect 1794 291454 2414 326898
rect 1794 290898 1826 291454
rect 2382 290898 2414 291454
rect 1794 255454 2414 290898
rect 1794 254898 1826 255454
rect 2382 254898 2414 255454
rect 1794 219454 2414 254898
rect 1794 218898 1826 219454
rect 2382 218898 2414 219454
rect 1794 183454 2414 218898
rect 1794 182898 1826 183454
rect 2382 182898 2414 183454
rect 1794 147454 2414 182898
rect 1794 146898 1826 147454
rect 2382 146898 2414 147454
rect 1794 111454 2414 146898
rect 1794 110898 1826 111454
rect 2382 110898 2414 111454
rect 1794 75454 2414 110898
rect 1794 74898 1826 75454
rect 2382 74898 2414 75454
rect 1794 39454 2414 74898
rect 1794 38898 1826 39454
rect 2382 38898 2414 39454
rect 1794 3454 2414 38898
rect 1794 2898 1826 3454
rect 2382 2898 2414 3454
rect 1794 -346 2414 2898
rect 1794 -902 1826 -346
rect 2382 -902 2414 -346
rect -2966 -1862 -2934 -1306
rect -2378 -1862 -2346 -1306
rect -2966 -1894 -2346 -1862
rect 1794 -1894 2414 -902
rect 5514 691174 6134 706202
rect 5514 690618 5546 691174
rect 6102 690618 6134 691174
rect 5514 655174 6134 690618
rect 5514 654618 5546 655174
rect 6102 654618 6134 655174
rect 5514 619174 6134 654618
rect 5514 618618 5546 619174
rect 6102 618618 6134 619174
rect 5514 583174 6134 618618
rect 5514 582618 5546 583174
rect 6102 582618 6134 583174
rect 5514 547174 6134 582618
rect 5514 546618 5546 547174
rect 6102 546618 6134 547174
rect 5514 511174 6134 546618
rect 5514 510618 5546 511174
rect 6102 510618 6134 511174
rect 5514 475174 6134 510618
rect 5514 474618 5546 475174
rect 6102 474618 6134 475174
rect 5514 439174 6134 474618
rect 5514 438618 5546 439174
rect 6102 438618 6134 439174
rect 5514 403174 6134 438618
rect 5514 402618 5546 403174
rect 6102 402618 6134 403174
rect 5514 367174 6134 402618
rect 5514 366618 5546 367174
rect 6102 366618 6134 367174
rect 5514 331174 6134 366618
rect 5514 330618 5546 331174
rect 6102 330618 6134 331174
rect 5514 295174 6134 330618
rect 5514 294618 5546 295174
rect 6102 294618 6134 295174
rect 5514 259174 6134 294618
rect 5514 258618 5546 259174
rect 6102 258618 6134 259174
rect 5514 223174 6134 258618
rect 5514 222618 5546 223174
rect 6102 222618 6134 223174
rect 5514 187174 6134 222618
rect 5514 186618 5546 187174
rect 6102 186618 6134 187174
rect 5514 151174 6134 186618
rect 5514 150618 5546 151174
rect 6102 150618 6134 151174
rect 5514 115174 6134 150618
rect 5514 114618 5546 115174
rect 6102 114618 6134 115174
rect 5514 79174 6134 114618
rect 5514 78618 5546 79174
rect 6102 78618 6134 79174
rect 5514 43174 6134 78618
rect 5514 42618 5546 43174
rect 6102 42618 6134 43174
rect 5514 7174 6134 42618
rect 5514 6618 5546 7174
rect 6102 6618 6134 7174
rect -3926 -2822 -3894 -2266
rect -3338 -2822 -3306 -2266
rect -3926 -2854 -3306 -2822
rect 5514 -2266 6134 6618
rect 5514 -2822 5546 -2266
rect 6102 -2822 6134 -2266
rect -4886 -3782 -4854 -3226
rect -4298 -3782 -4266 -3226
rect -4886 -3814 -4266 -3782
rect 5514 -3814 6134 -2822
rect 9234 694894 9854 708122
rect 9234 694338 9266 694894
rect 9822 694338 9854 694894
rect 9234 658894 9854 694338
rect 9234 658338 9266 658894
rect 9822 658338 9854 658894
rect 9234 622894 9854 658338
rect 9234 622338 9266 622894
rect 9822 622338 9854 622894
rect 9234 586894 9854 622338
rect 9234 586338 9266 586894
rect 9822 586338 9854 586894
rect 9234 550894 9854 586338
rect 9234 550338 9266 550894
rect 9822 550338 9854 550894
rect 9234 514894 9854 550338
rect 9234 514338 9266 514894
rect 9822 514338 9854 514894
rect 9234 478894 9854 514338
rect 9234 478338 9266 478894
rect 9822 478338 9854 478894
rect 9234 442894 9854 478338
rect 9234 442338 9266 442894
rect 9822 442338 9854 442894
rect 9234 406894 9854 442338
rect 9234 406338 9266 406894
rect 9822 406338 9854 406894
rect 9234 370894 9854 406338
rect 9234 370338 9266 370894
rect 9822 370338 9854 370894
rect 9234 334894 9854 370338
rect 9234 334338 9266 334894
rect 9822 334338 9854 334894
rect 9234 298894 9854 334338
rect 9234 298338 9266 298894
rect 9822 298338 9854 298894
rect 9234 262894 9854 298338
rect 9234 262338 9266 262894
rect 9822 262338 9854 262894
rect 9234 226894 9854 262338
rect 9234 226338 9266 226894
rect 9822 226338 9854 226894
rect 9234 190894 9854 226338
rect 9234 190338 9266 190894
rect 9822 190338 9854 190894
rect 9234 154894 9854 190338
rect 9234 154338 9266 154894
rect 9822 154338 9854 154894
rect 9234 118894 9854 154338
rect 9234 118338 9266 118894
rect 9822 118338 9854 118894
rect 9234 82894 9854 118338
rect 9234 82338 9266 82894
rect 9822 82338 9854 82894
rect 9234 46894 9854 82338
rect 9234 46338 9266 46894
rect 9822 46338 9854 46894
rect 9234 10894 9854 46338
rect 9234 10338 9266 10894
rect 9822 10338 9854 10894
rect -5846 -4742 -5814 -4186
rect -5258 -4742 -5226 -4186
rect -5846 -4774 -5226 -4742
rect 9234 -4186 9854 10338
rect 9234 -4742 9266 -4186
rect 9822 -4742 9854 -4186
rect -6806 -5702 -6774 -5146
rect -6218 -5702 -6186 -5146
rect -6806 -5734 -6186 -5702
rect 9234 -5734 9854 -4742
rect 12954 698614 13574 710042
rect 30954 711558 31574 711590
rect 30954 711002 30986 711558
rect 31542 711002 31574 711558
rect 27234 709638 27854 709670
rect 27234 709082 27266 709638
rect 27822 709082 27854 709638
rect 23514 707718 24134 707750
rect 23514 707162 23546 707718
rect 24102 707162 24134 707718
rect 12954 698058 12986 698614
rect 13542 698058 13574 698614
rect 12954 662614 13574 698058
rect 12954 662058 12986 662614
rect 13542 662058 13574 662614
rect 12954 626614 13574 662058
rect 12954 626058 12986 626614
rect 13542 626058 13574 626614
rect 12954 590614 13574 626058
rect 12954 590058 12986 590614
rect 13542 590058 13574 590614
rect 12954 554614 13574 590058
rect 12954 554058 12986 554614
rect 13542 554058 13574 554614
rect 12954 518614 13574 554058
rect 12954 518058 12986 518614
rect 13542 518058 13574 518614
rect 12954 482614 13574 518058
rect 12954 482058 12986 482614
rect 13542 482058 13574 482614
rect 12954 446614 13574 482058
rect 12954 446058 12986 446614
rect 13542 446058 13574 446614
rect 12954 410614 13574 446058
rect 12954 410058 12986 410614
rect 13542 410058 13574 410614
rect 12954 374614 13574 410058
rect 12954 374058 12986 374614
rect 13542 374058 13574 374614
rect 12954 338614 13574 374058
rect 12954 338058 12986 338614
rect 13542 338058 13574 338614
rect 12954 302614 13574 338058
rect 12954 302058 12986 302614
rect 13542 302058 13574 302614
rect 12954 266614 13574 302058
rect 12954 266058 12986 266614
rect 13542 266058 13574 266614
rect 12954 230614 13574 266058
rect 12954 230058 12986 230614
rect 13542 230058 13574 230614
rect 12954 194614 13574 230058
rect 12954 194058 12986 194614
rect 13542 194058 13574 194614
rect 12954 158614 13574 194058
rect 12954 158058 12986 158614
rect 13542 158058 13574 158614
rect 12954 122614 13574 158058
rect 12954 122058 12986 122614
rect 13542 122058 13574 122614
rect 12954 86614 13574 122058
rect 12954 86058 12986 86614
rect 13542 86058 13574 86614
rect 12954 50614 13574 86058
rect 12954 50058 12986 50614
rect 13542 50058 13574 50614
rect 12954 14614 13574 50058
rect 12954 14058 12986 14614
rect 13542 14058 13574 14614
rect -7766 -6662 -7734 -6106
rect -7178 -6662 -7146 -6106
rect -7766 -6694 -7146 -6662
rect 12954 -6106 13574 14058
rect 19794 705798 20414 705830
rect 19794 705242 19826 705798
rect 20382 705242 20414 705798
rect 19794 669454 20414 705242
rect 19794 668898 19826 669454
rect 20382 668898 20414 669454
rect 19794 633454 20414 668898
rect 19794 632898 19826 633454
rect 20382 632898 20414 633454
rect 19794 597454 20414 632898
rect 19794 596898 19826 597454
rect 20382 596898 20414 597454
rect 19794 561454 20414 596898
rect 19794 560898 19826 561454
rect 20382 560898 20414 561454
rect 19794 525454 20414 560898
rect 19794 524898 19826 525454
rect 20382 524898 20414 525454
rect 19794 489454 20414 524898
rect 19794 488898 19826 489454
rect 20382 488898 20414 489454
rect 19794 453454 20414 488898
rect 19794 452898 19826 453454
rect 20382 452898 20414 453454
rect 19794 417454 20414 452898
rect 19794 416898 19826 417454
rect 20382 416898 20414 417454
rect 19794 381454 20414 416898
rect 19794 380898 19826 381454
rect 20382 380898 20414 381454
rect 19794 345454 20414 380898
rect 19794 344898 19826 345454
rect 20382 344898 20414 345454
rect 19794 309454 20414 344898
rect 19794 308898 19826 309454
rect 20382 308898 20414 309454
rect 19794 273454 20414 308898
rect 19794 272898 19826 273454
rect 20382 272898 20414 273454
rect 19794 237454 20414 272898
rect 19794 236898 19826 237454
rect 20382 236898 20414 237454
rect 19794 201454 20414 236898
rect 19794 200898 19826 201454
rect 20382 200898 20414 201454
rect 19794 165454 20414 200898
rect 19794 164898 19826 165454
rect 20382 164898 20414 165454
rect 19794 129454 20414 164898
rect 19794 128898 19826 129454
rect 20382 128898 20414 129454
rect 19794 93454 20414 128898
rect 19794 92898 19826 93454
rect 20382 92898 20414 93454
rect 19794 57454 20414 92898
rect 19794 56898 19826 57454
rect 20382 56898 20414 57454
rect 19794 21454 20414 56898
rect 19794 20898 19826 21454
rect 20382 20898 20414 21454
rect 19794 -1306 20414 20898
rect 19794 -1862 19826 -1306
rect 20382 -1862 20414 -1306
rect 19794 -1894 20414 -1862
rect 23514 673174 24134 707162
rect 23514 672618 23546 673174
rect 24102 672618 24134 673174
rect 23514 637174 24134 672618
rect 23514 636618 23546 637174
rect 24102 636618 24134 637174
rect 23514 601174 24134 636618
rect 23514 600618 23546 601174
rect 24102 600618 24134 601174
rect 23514 565174 24134 600618
rect 23514 564618 23546 565174
rect 24102 564618 24134 565174
rect 23514 529174 24134 564618
rect 23514 528618 23546 529174
rect 24102 528618 24134 529174
rect 23514 493174 24134 528618
rect 23514 492618 23546 493174
rect 24102 492618 24134 493174
rect 23514 457174 24134 492618
rect 23514 456618 23546 457174
rect 24102 456618 24134 457174
rect 23514 421174 24134 456618
rect 23514 420618 23546 421174
rect 24102 420618 24134 421174
rect 23514 385174 24134 420618
rect 23514 384618 23546 385174
rect 24102 384618 24134 385174
rect 23514 349174 24134 384618
rect 23514 348618 23546 349174
rect 24102 348618 24134 349174
rect 23514 313174 24134 348618
rect 23514 312618 23546 313174
rect 24102 312618 24134 313174
rect 23514 277174 24134 312618
rect 23514 276618 23546 277174
rect 24102 276618 24134 277174
rect 23514 241174 24134 276618
rect 23514 240618 23546 241174
rect 24102 240618 24134 241174
rect 23514 205174 24134 240618
rect 23514 204618 23546 205174
rect 24102 204618 24134 205174
rect 23514 169174 24134 204618
rect 23514 168618 23546 169174
rect 24102 168618 24134 169174
rect 23514 133174 24134 168618
rect 23514 132618 23546 133174
rect 24102 132618 24134 133174
rect 23514 97174 24134 132618
rect 23514 96618 23546 97174
rect 24102 96618 24134 97174
rect 23514 61174 24134 96618
rect 23514 60618 23546 61174
rect 24102 60618 24134 61174
rect 23514 25174 24134 60618
rect 23514 24618 23546 25174
rect 24102 24618 24134 25174
rect 23514 -3226 24134 24618
rect 23514 -3782 23546 -3226
rect 24102 -3782 24134 -3226
rect 23514 -3814 24134 -3782
rect 27234 676894 27854 709082
rect 27234 676338 27266 676894
rect 27822 676338 27854 676894
rect 27234 640894 27854 676338
rect 27234 640338 27266 640894
rect 27822 640338 27854 640894
rect 27234 604894 27854 640338
rect 27234 604338 27266 604894
rect 27822 604338 27854 604894
rect 27234 568894 27854 604338
rect 27234 568338 27266 568894
rect 27822 568338 27854 568894
rect 27234 532894 27854 568338
rect 27234 532338 27266 532894
rect 27822 532338 27854 532894
rect 27234 496894 27854 532338
rect 27234 496338 27266 496894
rect 27822 496338 27854 496894
rect 27234 460894 27854 496338
rect 27234 460338 27266 460894
rect 27822 460338 27854 460894
rect 27234 424894 27854 460338
rect 27234 424338 27266 424894
rect 27822 424338 27854 424894
rect 27234 388894 27854 424338
rect 27234 388338 27266 388894
rect 27822 388338 27854 388894
rect 27234 352894 27854 388338
rect 27234 352338 27266 352894
rect 27822 352338 27854 352894
rect 27234 316894 27854 352338
rect 27234 316338 27266 316894
rect 27822 316338 27854 316894
rect 27234 280894 27854 316338
rect 27234 280338 27266 280894
rect 27822 280338 27854 280894
rect 27234 244894 27854 280338
rect 27234 244338 27266 244894
rect 27822 244338 27854 244894
rect 27234 208894 27854 244338
rect 27234 208338 27266 208894
rect 27822 208338 27854 208894
rect 27234 172894 27854 208338
rect 27234 172338 27266 172894
rect 27822 172338 27854 172894
rect 27234 136894 27854 172338
rect 27234 136338 27266 136894
rect 27822 136338 27854 136894
rect 27234 100894 27854 136338
rect 27234 100338 27266 100894
rect 27822 100338 27854 100894
rect 27234 64894 27854 100338
rect 27234 64338 27266 64894
rect 27822 64338 27854 64894
rect 27234 28894 27854 64338
rect 27234 28338 27266 28894
rect 27822 28338 27854 28894
rect 27234 -5146 27854 28338
rect 27234 -5702 27266 -5146
rect 27822 -5702 27854 -5146
rect 27234 -5734 27854 -5702
rect 30954 680614 31574 711002
rect 48954 710598 49574 711590
rect 48954 710042 48986 710598
rect 49542 710042 49574 710598
rect 45234 708678 45854 709670
rect 45234 708122 45266 708678
rect 45822 708122 45854 708678
rect 41514 706758 42134 707750
rect 41514 706202 41546 706758
rect 42102 706202 42134 706758
rect 30954 680058 30986 680614
rect 31542 680058 31574 680614
rect 30954 644614 31574 680058
rect 30954 644058 30986 644614
rect 31542 644058 31574 644614
rect 30954 608614 31574 644058
rect 30954 608058 30986 608614
rect 31542 608058 31574 608614
rect 30954 572614 31574 608058
rect 30954 572058 30986 572614
rect 31542 572058 31574 572614
rect 30954 536614 31574 572058
rect 30954 536058 30986 536614
rect 31542 536058 31574 536614
rect 30954 500614 31574 536058
rect 30954 500058 30986 500614
rect 31542 500058 31574 500614
rect 30954 464614 31574 500058
rect 30954 464058 30986 464614
rect 31542 464058 31574 464614
rect 30954 428614 31574 464058
rect 30954 428058 30986 428614
rect 31542 428058 31574 428614
rect 30954 392614 31574 428058
rect 30954 392058 30986 392614
rect 31542 392058 31574 392614
rect 30954 356614 31574 392058
rect 30954 356058 30986 356614
rect 31542 356058 31574 356614
rect 30954 320614 31574 356058
rect 30954 320058 30986 320614
rect 31542 320058 31574 320614
rect 30954 284614 31574 320058
rect 30954 284058 30986 284614
rect 31542 284058 31574 284614
rect 30954 248614 31574 284058
rect 30954 248058 30986 248614
rect 31542 248058 31574 248614
rect 30954 212614 31574 248058
rect 30954 212058 30986 212614
rect 31542 212058 31574 212614
rect 30954 176614 31574 212058
rect 30954 176058 30986 176614
rect 31542 176058 31574 176614
rect 30954 140614 31574 176058
rect 30954 140058 30986 140614
rect 31542 140058 31574 140614
rect 30954 104614 31574 140058
rect 30954 104058 30986 104614
rect 31542 104058 31574 104614
rect 30954 68614 31574 104058
rect 30954 68058 30986 68614
rect 31542 68058 31574 68614
rect 30954 32614 31574 68058
rect 30954 32058 30986 32614
rect 31542 32058 31574 32614
rect 12954 -6662 12986 -6106
rect 13542 -6662 13574 -6106
rect -8726 -7622 -8694 -7066
rect -8138 -7622 -8106 -7066
rect -8726 -7654 -8106 -7622
rect 12954 -7654 13574 -6662
rect 30954 -7066 31574 32058
rect 37794 704838 38414 705830
rect 37794 704282 37826 704838
rect 38382 704282 38414 704838
rect 37794 687454 38414 704282
rect 37794 686898 37826 687454
rect 38382 686898 38414 687454
rect 37794 651454 38414 686898
rect 37794 650898 37826 651454
rect 38382 650898 38414 651454
rect 37794 615454 38414 650898
rect 37794 614898 37826 615454
rect 38382 614898 38414 615454
rect 37794 579454 38414 614898
rect 37794 578898 37826 579454
rect 38382 578898 38414 579454
rect 37794 543454 38414 578898
rect 37794 542898 37826 543454
rect 38382 542898 38414 543454
rect 37794 507454 38414 542898
rect 37794 506898 37826 507454
rect 38382 506898 38414 507454
rect 37794 471454 38414 506898
rect 37794 470898 37826 471454
rect 38382 470898 38414 471454
rect 37794 435454 38414 470898
rect 37794 434898 37826 435454
rect 38382 434898 38414 435454
rect 37794 399454 38414 434898
rect 37794 398898 37826 399454
rect 38382 398898 38414 399454
rect 37794 363454 38414 398898
rect 37794 362898 37826 363454
rect 38382 362898 38414 363454
rect 37794 327454 38414 362898
rect 37794 326898 37826 327454
rect 38382 326898 38414 327454
rect 37794 291454 38414 326898
rect 37794 290898 37826 291454
rect 38382 290898 38414 291454
rect 37794 255454 38414 290898
rect 37794 254898 37826 255454
rect 38382 254898 38414 255454
rect 37794 219454 38414 254898
rect 37794 218898 37826 219454
rect 38382 218898 38414 219454
rect 37794 183454 38414 218898
rect 37794 182898 37826 183454
rect 38382 182898 38414 183454
rect 37794 147454 38414 182898
rect 37794 146898 37826 147454
rect 38382 146898 38414 147454
rect 37794 111454 38414 146898
rect 37794 110898 37826 111454
rect 38382 110898 38414 111454
rect 37794 75454 38414 110898
rect 37794 74898 37826 75454
rect 38382 74898 38414 75454
rect 37794 39454 38414 74898
rect 37794 38898 37826 39454
rect 38382 38898 38414 39454
rect 37794 3454 38414 38898
rect 37794 2898 37826 3454
rect 38382 2898 38414 3454
rect 37794 -346 38414 2898
rect 37794 -902 37826 -346
rect 38382 -902 38414 -346
rect 37794 -1894 38414 -902
rect 41514 691174 42134 706202
rect 41514 690618 41546 691174
rect 42102 690618 42134 691174
rect 41514 655174 42134 690618
rect 41514 654618 41546 655174
rect 42102 654618 42134 655174
rect 41514 619174 42134 654618
rect 41514 618618 41546 619174
rect 42102 618618 42134 619174
rect 41514 583174 42134 618618
rect 41514 582618 41546 583174
rect 42102 582618 42134 583174
rect 41514 547174 42134 582618
rect 41514 546618 41546 547174
rect 42102 546618 42134 547174
rect 41514 511174 42134 546618
rect 41514 510618 41546 511174
rect 42102 510618 42134 511174
rect 41514 475174 42134 510618
rect 41514 474618 41546 475174
rect 42102 474618 42134 475174
rect 41514 439174 42134 474618
rect 41514 438618 41546 439174
rect 42102 438618 42134 439174
rect 41514 403174 42134 438618
rect 41514 402618 41546 403174
rect 42102 402618 42134 403174
rect 41514 367174 42134 402618
rect 41514 366618 41546 367174
rect 42102 366618 42134 367174
rect 41514 331174 42134 366618
rect 41514 330618 41546 331174
rect 42102 330618 42134 331174
rect 41514 295174 42134 330618
rect 41514 294618 41546 295174
rect 42102 294618 42134 295174
rect 41514 259174 42134 294618
rect 41514 258618 41546 259174
rect 42102 258618 42134 259174
rect 41514 223174 42134 258618
rect 41514 222618 41546 223174
rect 42102 222618 42134 223174
rect 41514 187174 42134 222618
rect 41514 186618 41546 187174
rect 42102 186618 42134 187174
rect 41514 151174 42134 186618
rect 41514 150618 41546 151174
rect 42102 150618 42134 151174
rect 41514 115174 42134 150618
rect 41514 114618 41546 115174
rect 42102 114618 42134 115174
rect 41514 79174 42134 114618
rect 41514 78618 41546 79174
rect 42102 78618 42134 79174
rect 41514 43174 42134 78618
rect 41514 42618 41546 43174
rect 42102 42618 42134 43174
rect 41514 7174 42134 42618
rect 41514 6618 41546 7174
rect 42102 6618 42134 7174
rect 41514 -2266 42134 6618
rect 41514 -2822 41546 -2266
rect 42102 -2822 42134 -2266
rect 41514 -3814 42134 -2822
rect 45234 694894 45854 708122
rect 45234 694338 45266 694894
rect 45822 694338 45854 694894
rect 45234 658894 45854 694338
rect 45234 658338 45266 658894
rect 45822 658338 45854 658894
rect 45234 622894 45854 658338
rect 45234 622338 45266 622894
rect 45822 622338 45854 622894
rect 45234 586894 45854 622338
rect 45234 586338 45266 586894
rect 45822 586338 45854 586894
rect 45234 550894 45854 586338
rect 45234 550338 45266 550894
rect 45822 550338 45854 550894
rect 45234 514894 45854 550338
rect 45234 514338 45266 514894
rect 45822 514338 45854 514894
rect 45234 478894 45854 514338
rect 45234 478338 45266 478894
rect 45822 478338 45854 478894
rect 45234 442894 45854 478338
rect 45234 442338 45266 442894
rect 45822 442338 45854 442894
rect 45234 406894 45854 442338
rect 45234 406338 45266 406894
rect 45822 406338 45854 406894
rect 45234 370894 45854 406338
rect 45234 370338 45266 370894
rect 45822 370338 45854 370894
rect 45234 334894 45854 370338
rect 45234 334338 45266 334894
rect 45822 334338 45854 334894
rect 45234 298894 45854 334338
rect 45234 298338 45266 298894
rect 45822 298338 45854 298894
rect 45234 262894 45854 298338
rect 45234 262338 45266 262894
rect 45822 262338 45854 262894
rect 45234 226894 45854 262338
rect 45234 226338 45266 226894
rect 45822 226338 45854 226894
rect 45234 190894 45854 226338
rect 45234 190338 45266 190894
rect 45822 190338 45854 190894
rect 45234 154894 45854 190338
rect 45234 154338 45266 154894
rect 45822 154338 45854 154894
rect 45234 118894 45854 154338
rect 45234 118338 45266 118894
rect 45822 118338 45854 118894
rect 45234 82894 45854 118338
rect 45234 82338 45266 82894
rect 45822 82338 45854 82894
rect 45234 46894 45854 82338
rect 45234 46338 45266 46894
rect 45822 46338 45854 46894
rect 45234 10894 45854 46338
rect 45234 10338 45266 10894
rect 45822 10338 45854 10894
rect 45234 -4186 45854 10338
rect 45234 -4742 45266 -4186
rect 45822 -4742 45854 -4186
rect 45234 -5734 45854 -4742
rect 48954 698614 49574 710042
rect 66954 711558 67574 711590
rect 66954 711002 66986 711558
rect 67542 711002 67574 711558
rect 63234 709638 63854 709670
rect 63234 709082 63266 709638
rect 63822 709082 63854 709638
rect 59514 707718 60134 707750
rect 59514 707162 59546 707718
rect 60102 707162 60134 707718
rect 48954 698058 48986 698614
rect 49542 698058 49574 698614
rect 48954 662614 49574 698058
rect 48954 662058 48986 662614
rect 49542 662058 49574 662614
rect 48954 626614 49574 662058
rect 48954 626058 48986 626614
rect 49542 626058 49574 626614
rect 48954 590614 49574 626058
rect 48954 590058 48986 590614
rect 49542 590058 49574 590614
rect 48954 554614 49574 590058
rect 48954 554058 48986 554614
rect 49542 554058 49574 554614
rect 48954 518614 49574 554058
rect 48954 518058 48986 518614
rect 49542 518058 49574 518614
rect 48954 482614 49574 518058
rect 48954 482058 48986 482614
rect 49542 482058 49574 482614
rect 48954 446614 49574 482058
rect 48954 446058 48986 446614
rect 49542 446058 49574 446614
rect 48954 410614 49574 446058
rect 48954 410058 48986 410614
rect 49542 410058 49574 410614
rect 48954 374614 49574 410058
rect 48954 374058 48986 374614
rect 49542 374058 49574 374614
rect 48954 338614 49574 374058
rect 48954 338058 48986 338614
rect 49542 338058 49574 338614
rect 48954 302614 49574 338058
rect 48954 302058 48986 302614
rect 49542 302058 49574 302614
rect 48954 266614 49574 302058
rect 48954 266058 48986 266614
rect 49542 266058 49574 266614
rect 48954 230614 49574 266058
rect 48954 230058 48986 230614
rect 49542 230058 49574 230614
rect 48954 194614 49574 230058
rect 48954 194058 48986 194614
rect 49542 194058 49574 194614
rect 48954 158614 49574 194058
rect 48954 158058 48986 158614
rect 49542 158058 49574 158614
rect 48954 122614 49574 158058
rect 48954 122058 48986 122614
rect 49542 122058 49574 122614
rect 48954 86614 49574 122058
rect 48954 86058 48986 86614
rect 49542 86058 49574 86614
rect 48954 50614 49574 86058
rect 48954 50058 48986 50614
rect 49542 50058 49574 50614
rect 48954 14614 49574 50058
rect 48954 14058 48986 14614
rect 49542 14058 49574 14614
rect 30954 -7622 30986 -7066
rect 31542 -7622 31574 -7066
rect 30954 -7654 31574 -7622
rect 48954 -6106 49574 14058
rect 55794 705798 56414 705830
rect 55794 705242 55826 705798
rect 56382 705242 56414 705798
rect 55794 669454 56414 705242
rect 55794 668898 55826 669454
rect 56382 668898 56414 669454
rect 55794 633454 56414 668898
rect 55794 632898 55826 633454
rect 56382 632898 56414 633454
rect 55794 597454 56414 632898
rect 55794 596898 55826 597454
rect 56382 596898 56414 597454
rect 55794 561454 56414 596898
rect 55794 560898 55826 561454
rect 56382 560898 56414 561454
rect 55794 525454 56414 560898
rect 55794 524898 55826 525454
rect 56382 524898 56414 525454
rect 55794 489454 56414 524898
rect 55794 488898 55826 489454
rect 56382 488898 56414 489454
rect 55794 453454 56414 488898
rect 55794 452898 55826 453454
rect 56382 452898 56414 453454
rect 55794 417454 56414 452898
rect 55794 416898 55826 417454
rect 56382 416898 56414 417454
rect 55794 381454 56414 416898
rect 55794 380898 55826 381454
rect 56382 380898 56414 381454
rect 55794 345454 56414 380898
rect 55794 344898 55826 345454
rect 56382 344898 56414 345454
rect 55794 309454 56414 344898
rect 55794 308898 55826 309454
rect 56382 308898 56414 309454
rect 55794 273454 56414 308898
rect 55794 272898 55826 273454
rect 56382 272898 56414 273454
rect 55794 237454 56414 272898
rect 55794 236898 55826 237454
rect 56382 236898 56414 237454
rect 55794 201454 56414 236898
rect 55794 200898 55826 201454
rect 56382 200898 56414 201454
rect 55794 165454 56414 200898
rect 55794 164898 55826 165454
rect 56382 164898 56414 165454
rect 55794 129454 56414 164898
rect 55794 128898 55826 129454
rect 56382 128898 56414 129454
rect 55794 93454 56414 128898
rect 55794 92898 55826 93454
rect 56382 92898 56414 93454
rect 55794 57454 56414 92898
rect 55794 56898 55826 57454
rect 56382 56898 56414 57454
rect 55794 21454 56414 56898
rect 55794 20898 55826 21454
rect 56382 20898 56414 21454
rect 55794 -1306 56414 20898
rect 55794 -1862 55826 -1306
rect 56382 -1862 56414 -1306
rect 55794 -1894 56414 -1862
rect 59514 673174 60134 707162
rect 59514 672618 59546 673174
rect 60102 672618 60134 673174
rect 59514 637174 60134 672618
rect 59514 636618 59546 637174
rect 60102 636618 60134 637174
rect 59514 601174 60134 636618
rect 59514 600618 59546 601174
rect 60102 600618 60134 601174
rect 59514 565174 60134 600618
rect 59514 564618 59546 565174
rect 60102 564618 60134 565174
rect 59514 529174 60134 564618
rect 59514 528618 59546 529174
rect 60102 528618 60134 529174
rect 59514 493174 60134 528618
rect 59514 492618 59546 493174
rect 60102 492618 60134 493174
rect 59514 457174 60134 492618
rect 59514 456618 59546 457174
rect 60102 456618 60134 457174
rect 59514 421174 60134 456618
rect 59514 420618 59546 421174
rect 60102 420618 60134 421174
rect 59514 385174 60134 420618
rect 59514 384618 59546 385174
rect 60102 384618 60134 385174
rect 59514 349174 60134 384618
rect 59514 348618 59546 349174
rect 60102 348618 60134 349174
rect 59514 313174 60134 348618
rect 59514 312618 59546 313174
rect 60102 312618 60134 313174
rect 59514 277174 60134 312618
rect 59514 276618 59546 277174
rect 60102 276618 60134 277174
rect 59514 241174 60134 276618
rect 59514 240618 59546 241174
rect 60102 240618 60134 241174
rect 59514 205174 60134 240618
rect 59514 204618 59546 205174
rect 60102 204618 60134 205174
rect 59514 169174 60134 204618
rect 59514 168618 59546 169174
rect 60102 168618 60134 169174
rect 59514 133174 60134 168618
rect 59514 132618 59546 133174
rect 60102 132618 60134 133174
rect 59514 97174 60134 132618
rect 59514 96618 59546 97174
rect 60102 96618 60134 97174
rect 59514 61174 60134 96618
rect 59514 60618 59546 61174
rect 60102 60618 60134 61174
rect 59514 25174 60134 60618
rect 59514 24618 59546 25174
rect 60102 24618 60134 25174
rect 59514 -3226 60134 24618
rect 59514 -3782 59546 -3226
rect 60102 -3782 60134 -3226
rect 59514 -3814 60134 -3782
rect 63234 676894 63854 709082
rect 63234 676338 63266 676894
rect 63822 676338 63854 676894
rect 63234 640894 63854 676338
rect 63234 640338 63266 640894
rect 63822 640338 63854 640894
rect 63234 604894 63854 640338
rect 63234 604338 63266 604894
rect 63822 604338 63854 604894
rect 63234 568894 63854 604338
rect 63234 568338 63266 568894
rect 63822 568338 63854 568894
rect 63234 532894 63854 568338
rect 63234 532338 63266 532894
rect 63822 532338 63854 532894
rect 63234 496894 63854 532338
rect 63234 496338 63266 496894
rect 63822 496338 63854 496894
rect 63234 460894 63854 496338
rect 63234 460338 63266 460894
rect 63822 460338 63854 460894
rect 63234 424894 63854 460338
rect 63234 424338 63266 424894
rect 63822 424338 63854 424894
rect 63234 388894 63854 424338
rect 63234 388338 63266 388894
rect 63822 388338 63854 388894
rect 63234 352894 63854 388338
rect 63234 352338 63266 352894
rect 63822 352338 63854 352894
rect 63234 316894 63854 352338
rect 63234 316338 63266 316894
rect 63822 316338 63854 316894
rect 63234 280894 63854 316338
rect 63234 280338 63266 280894
rect 63822 280338 63854 280894
rect 63234 244894 63854 280338
rect 63234 244338 63266 244894
rect 63822 244338 63854 244894
rect 63234 208894 63854 244338
rect 63234 208338 63266 208894
rect 63822 208338 63854 208894
rect 63234 172894 63854 208338
rect 63234 172338 63266 172894
rect 63822 172338 63854 172894
rect 63234 136894 63854 172338
rect 63234 136338 63266 136894
rect 63822 136338 63854 136894
rect 63234 100894 63854 136338
rect 63234 100338 63266 100894
rect 63822 100338 63854 100894
rect 63234 64894 63854 100338
rect 63234 64338 63266 64894
rect 63822 64338 63854 64894
rect 63234 28894 63854 64338
rect 63234 28338 63266 28894
rect 63822 28338 63854 28894
rect 63234 -5146 63854 28338
rect 63234 -5702 63266 -5146
rect 63822 -5702 63854 -5146
rect 63234 -5734 63854 -5702
rect 66954 680614 67574 711002
rect 84954 710598 85574 711590
rect 84954 710042 84986 710598
rect 85542 710042 85574 710598
rect 81234 708678 81854 709670
rect 81234 708122 81266 708678
rect 81822 708122 81854 708678
rect 77514 706758 78134 707750
rect 77514 706202 77546 706758
rect 78102 706202 78134 706758
rect 66954 680058 66986 680614
rect 67542 680058 67574 680614
rect 66954 644614 67574 680058
rect 66954 644058 66986 644614
rect 67542 644058 67574 644614
rect 66954 608614 67574 644058
rect 66954 608058 66986 608614
rect 67542 608058 67574 608614
rect 66954 572614 67574 608058
rect 66954 572058 66986 572614
rect 67542 572058 67574 572614
rect 66954 536614 67574 572058
rect 66954 536058 66986 536614
rect 67542 536058 67574 536614
rect 66954 500614 67574 536058
rect 66954 500058 66986 500614
rect 67542 500058 67574 500614
rect 66954 464614 67574 500058
rect 66954 464058 66986 464614
rect 67542 464058 67574 464614
rect 66954 428614 67574 464058
rect 66954 428058 66986 428614
rect 67542 428058 67574 428614
rect 66954 392614 67574 428058
rect 66954 392058 66986 392614
rect 67542 392058 67574 392614
rect 66954 356614 67574 392058
rect 66954 356058 66986 356614
rect 67542 356058 67574 356614
rect 66954 320614 67574 356058
rect 66954 320058 66986 320614
rect 67542 320058 67574 320614
rect 66954 284614 67574 320058
rect 66954 284058 66986 284614
rect 67542 284058 67574 284614
rect 66954 248614 67574 284058
rect 66954 248058 66986 248614
rect 67542 248058 67574 248614
rect 66954 212614 67574 248058
rect 66954 212058 66986 212614
rect 67542 212058 67574 212614
rect 66954 176614 67574 212058
rect 66954 176058 66986 176614
rect 67542 176058 67574 176614
rect 66954 140614 67574 176058
rect 66954 140058 66986 140614
rect 67542 140058 67574 140614
rect 66954 104614 67574 140058
rect 66954 104058 66986 104614
rect 67542 104058 67574 104614
rect 66954 68614 67574 104058
rect 66954 68058 66986 68614
rect 67542 68058 67574 68614
rect 66954 32614 67574 68058
rect 66954 32058 66986 32614
rect 67542 32058 67574 32614
rect 48954 -6662 48986 -6106
rect 49542 -6662 49574 -6106
rect 48954 -7654 49574 -6662
rect 66954 -7066 67574 32058
rect 73794 704838 74414 705830
rect 73794 704282 73826 704838
rect 74382 704282 74414 704838
rect 73794 687454 74414 704282
rect 73794 686898 73826 687454
rect 74382 686898 74414 687454
rect 73794 651454 74414 686898
rect 73794 650898 73826 651454
rect 74382 650898 74414 651454
rect 73794 615454 74414 650898
rect 73794 614898 73826 615454
rect 74382 614898 74414 615454
rect 73794 579454 74414 614898
rect 73794 578898 73826 579454
rect 74382 578898 74414 579454
rect 73794 543454 74414 578898
rect 73794 542898 73826 543454
rect 74382 542898 74414 543454
rect 73794 507454 74414 542898
rect 73794 506898 73826 507454
rect 74382 506898 74414 507454
rect 73794 471454 74414 506898
rect 73794 470898 73826 471454
rect 74382 470898 74414 471454
rect 73794 435454 74414 470898
rect 73794 434898 73826 435454
rect 74382 434898 74414 435454
rect 73794 399454 74414 434898
rect 73794 398898 73826 399454
rect 74382 398898 74414 399454
rect 73794 363454 74414 398898
rect 73794 362898 73826 363454
rect 74382 362898 74414 363454
rect 73794 327454 74414 362898
rect 73794 326898 73826 327454
rect 74382 326898 74414 327454
rect 73794 291454 74414 326898
rect 73794 290898 73826 291454
rect 74382 290898 74414 291454
rect 73794 255454 74414 290898
rect 73794 254898 73826 255454
rect 74382 254898 74414 255454
rect 73794 219454 74414 254898
rect 73794 218898 73826 219454
rect 74382 218898 74414 219454
rect 73794 183454 74414 218898
rect 73794 182898 73826 183454
rect 74382 182898 74414 183454
rect 73794 147454 74414 182898
rect 73794 146898 73826 147454
rect 74382 146898 74414 147454
rect 73794 111454 74414 146898
rect 73794 110898 73826 111454
rect 74382 110898 74414 111454
rect 73794 75454 74414 110898
rect 73794 74898 73826 75454
rect 74382 74898 74414 75454
rect 73794 39454 74414 74898
rect 73794 38898 73826 39454
rect 74382 38898 74414 39454
rect 73794 3454 74414 38898
rect 73794 2898 73826 3454
rect 74382 2898 74414 3454
rect 73794 -346 74414 2898
rect 73794 -902 73826 -346
rect 74382 -902 74414 -346
rect 73794 -1894 74414 -902
rect 77514 691174 78134 706202
rect 77514 690618 77546 691174
rect 78102 690618 78134 691174
rect 77514 655174 78134 690618
rect 77514 654618 77546 655174
rect 78102 654618 78134 655174
rect 77514 619174 78134 654618
rect 77514 618618 77546 619174
rect 78102 618618 78134 619174
rect 77514 583174 78134 618618
rect 77514 582618 77546 583174
rect 78102 582618 78134 583174
rect 77514 547174 78134 582618
rect 77514 546618 77546 547174
rect 78102 546618 78134 547174
rect 77514 511174 78134 546618
rect 77514 510618 77546 511174
rect 78102 510618 78134 511174
rect 77514 475174 78134 510618
rect 77514 474618 77546 475174
rect 78102 474618 78134 475174
rect 77514 439174 78134 474618
rect 77514 438618 77546 439174
rect 78102 438618 78134 439174
rect 77514 403174 78134 438618
rect 77514 402618 77546 403174
rect 78102 402618 78134 403174
rect 77514 367174 78134 402618
rect 77514 366618 77546 367174
rect 78102 366618 78134 367174
rect 77514 331174 78134 366618
rect 77514 330618 77546 331174
rect 78102 330618 78134 331174
rect 77514 295174 78134 330618
rect 77514 294618 77546 295174
rect 78102 294618 78134 295174
rect 77514 259174 78134 294618
rect 77514 258618 77546 259174
rect 78102 258618 78134 259174
rect 77514 223174 78134 258618
rect 77514 222618 77546 223174
rect 78102 222618 78134 223174
rect 77514 187174 78134 222618
rect 77514 186618 77546 187174
rect 78102 186618 78134 187174
rect 77514 151174 78134 186618
rect 77514 150618 77546 151174
rect 78102 150618 78134 151174
rect 77514 115174 78134 150618
rect 77514 114618 77546 115174
rect 78102 114618 78134 115174
rect 77514 79174 78134 114618
rect 77514 78618 77546 79174
rect 78102 78618 78134 79174
rect 77514 43174 78134 78618
rect 77514 42618 77546 43174
rect 78102 42618 78134 43174
rect 77514 7174 78134 42618
rect 77514 6618 77546 7174
rect 78102 6618 78134 7174
rect 77514 -2266 78134 6618
rect 77514 -2822 77546 -2266
rect 78102 -2822 78134 -2266
rect 77514 -3814 78134 -2822
rect 81234 694894 81854 708122
rect 81234 694338 81266 694894
rect 81822 694338 81854 694894
rect 81234 658894 81854 694338
rect 81234 658338 81266 658894
rect 81822 658338 81854 658894
rect 81234 622894 81854 658338
rect 81234 622338 81266 622894
rect 81822 622338 81854 622894
rect 81234 586894 81854 622338
rect 81234 586338 81266 586894
rect 81822 586338 81854 586894
rect 81234 550894 81854 586338
rect 81234 550338 81266 550894
rect 81822 550338 81854 550894
rect 81234 514894 81854 550338
rect 81234 514338 81266 514894
rect 81822 514338 81854 514894
rect 81234 478894 81854 514338
rect 81234 478338 81266 478894
rect 81822 478338 81854 478894
rect 81234 442894 81854 478338
rect 81234 442338 81266 442894
rect 81822 442338 81854 442894
rect 81234 406894 81854 442338
rect 81234 406338 81266 406894
rect 81822 406338 81854 406894
rect 81234 370894 81854 406338
rect 81234 370338 81266 370894
rect 81822 370338 81854 370894
rect 81234 334894 81854 370338
rect 81234 334338 81266 334894
rect 81822 334338 81854 334894
rect 81234 298894 81854 334338
rect 81234 298338 81266 298894
rect 81822 298338 81854 298894
rect 81234 262894 81854 298338
rect 81234 262338 81266 262894
rect 81822 262338 81854 262894
rect 81234 226894 81854 262338
rect 81234 226338 81266 226894
rect 81822 226338 81854 226894
rect 81234 190894 81854 226338
rect 81234 190338 81266 190894
rect 81822 190338 81854 190894
rect 81234 154894 81854 190338
rect 81234 154338 81266 154894
rect 81822 154338 81854 154894
rect 81234 118894 81854 154338
rect 81234 118338 81266 118894
rect 81822 118338 81854 118894
rect 81234 82894 81854 118338
rect 81234 82338 81266 82894
rect 81822 82338 81854 82894
rect 81234 46894 81854 82338
rect 81234 46338 81266 46894
rect 81822 46338 81854 46894
rect 81234 10894 81854 46338
rect 81234 10338 81266 10894
rect 81822 10338 81854 10894
rect 81234 -4186 81854 10338
rect 81234 -4742 81266 -4186
rect 81822 -4742 81854 -4186
rect 81234 -5734 81854 -4742
rect 84954 698614 85574 710042
rect 102954 711558 103574 711590
rect 102954 711002 102986 711558
rect 103542 711002 103574 711558
rect 99234 709638 99854 709670
rect 99234 709082 99266 709638
rect 99822 709082 99854 709638
rect 95514 707718 96134 707750
rect 95514 707162 95546 707718
rect 96102 707162 96134 707718
rect 84954 698058 84986 698614
rect 85542 698058 85574 698614
rect 84954 662614 85574 698058
rect 84954 662058 84986 662614
rect 85542 662058 85574 662614
rect 84954 626614 85574 662058
rect 84954 626058 84986 626614
rect 85542 626058 85574 626614
rect 84954 590614 85574 626058
rect 84954 590058 84986 590614
rect 85542 590058 85574 590614
rect 84954 554614 85574 590058
rect 84954 554058 84986 554614
rect 85542 554058 85574 554614
rect 84954 518614 85574 554058
rect 84954 518058 84986 518614
rect 85542 518058 85574 518614
rect 84954 482614 85574 518058
rect 84954 482058 84986 482614
rect 85542 482058 85574 482614
rect 84954 446614 85574 482058
rect 84954 446058 84986 446614
rect 85542 446058 85574 446614
rect 84954 410614 85574 446058
rect 84954 410058 84986 410614
rect 85542 410058 85574 410614
rect 84954 374614 85574 410058
rect 84954 374058 84986 374614
rect 85542 374058 85574 374614
rect 84954 338614 85574 374058
rect 84954 338058 84986 338614
rect 85542 338058 85574 338614
rect 84954 302614 85574 338058
rect 84954 302058 84986 302614
rect 85542 302058 85574 302614
rect 84954 266614 85574 302058
rect 84954 266058 84986 266614
rect 85542 266058 85574 266614
rect 84954 230614 85574 266058
rect 84954 230058 84986 230614
rect 85542 230058 85574 230614
rect 84954 194614 85574 230058
rect 84954 194058 84986 194614
rect 85542 194058 85574 194614
rect 84954 158614 85574 194058
rect 84954 158058 84986 158614
rect 85542 158058 85574 158614
rect 84954 122614 85574 158058
rect 84954 122058 84986 122614
rect 85542 122058 85574 122614
rect 84954 86614 85574 122058
rect 84954 86058 84986 86614
rect 85542 86058 85574 86614
rect 84954 50614 85574 86058
rect 84954 50058 84986 50614
rect 85542 50058 85574 50614
rect 84954 14614 85574 50058
rect 84954 14058 84986 14614
rect 85542 14058 85574 14614
rect 66954 -7622 66986 -7066
rect 67542 -7622 67574 -7066
rect 66954 -7654 67574 -7622
rect 84954 -6106 85574 14058
rect 91794 705798 92414 705830
rect 91794 705242 91826 705798
rect 92382 705242 92414 705798
rect 91794 669454 92414 705242
rect 91794 668898 91826 669454
rect 92382 668898 92414 669454
rect 91794 633454 92414 668898
rect 91794 632898 91826 633454
rect 92382 632898 92414 633454
rect 91794 597454 92414 632898
rect 91794 596898 91826 597454
rect 92382 596898 92414 597454
rect 91794 561454 92414 596898
rect 91794 560898 91826 561454
rect 92382 560898 92414 561454
rect 91794 525454 92414 560898
rect 91794 524898 91826 525454
rect 92382 524898 92414 525454
rect 91794 489454 92414 524898
rect 91794 488898 91826 489454
rect 92382 488898 92414 489454
rect 91794 453454 92414 488898
rect 91794 452898 91826 453454
rect 92382 452898 92414 453454
rect 91794 417454 92414 452898
rect 91794 416898 91826 417454
rect 92382 416898 92414 417454
rect 91794 381454 92414 416898
rect 91794 380898 91826 381454
rect 92382 380898 92414 381454
rect 91794 345454 92414 380898
rect 91794 344898 91826 345454
rect 92382 344898 92414 345454
rect 91794 309454 92414 344898
rect 91794 308898 91826 309454
rect 92382 308898 92414 309454
rect 91794 273454 92414 308898
rect 91794 272898 91826 273454
rect 92382 272898 92414 273454
rect 91794 237454 92414 272898
rect 91794 236898 91826 237454
rect 92382 236898 92414 237454
rect 91794 201454 92414 236898
rect 91794 200898 91826 201454
rect 92382 200898 92414 201454
rect 91794 165454 92414 200898
rect 91794 164898 91826 165454
rect 92382 164898 92414 165454
rect 91794 129454 92414 164898
rect 91794 128898 91826 129454
rect 92382 128898 92414 129454
rect 91794 93454 92414 128898
rect 91794 92898 91826 93454
rect 92382 92898 92414 93454
rect 91794 57454 92414 92898
rect 91794 56898 91826 57454
rect 92382 56898 92414 57454
rect 91794 21454 92414 56898
rect 91794 20898 91826 21454
rect 92382 20898 92414 21454
rect 91794 -1306 92414 20898
rect 91794 -1862 91826 -1306
rect 92382 -1862 92414 -1306
rect 91794 -1894 92414 -1862
rect 95514 673174 96134 707162
rect 95514 672618 95546 673174
rect 96102 672618 96134 673174
rect 95514 637174 96134 672618
rect 95514 636618 95546 637174
rect 96102 636618 96134 637174
rect 95514 601174 96134 636618
rect 95514 600618 95546 601174
rect 96102 600618 96134 601174
rect 95514 565174 96134 600618
rect 95514 564618 95546 565174
rect 96102 564618 96134 565174
rect 95514 529174 96134 564618
rect 95514 528618 95546 529174
rect 96102 528618 96134 529174
rect 95514 493174 96134 528618
rect 95514 492618 95546 493174
rect 96102 492618 96134 493174
rect 95514 457174 96134 492618
rect 95514 456618 95546 457174
rect 96102 456618 96134 457174
rect 95514 421174 96134 456618
rect 95514 420618 95546 421174
rect 96102 420618 96134 421174
rect 95514 385174 96134 420618
rect 95514 384618 95546 385174
rect 96102 384618 96134 385174
rect 95514 349174 96134 384618
rect 95514 348618 95546 349174
rect 96102 348618 96134 349174
rect 95514 313174 96134 348618
rect 95514 312618 95546 313174
rect 96102 312618 96134 313174
rect 95514 277174 96134 312618
rect 95514 276618 95546 277174
rect 96102 276618 96134 277174
rect 95514 241174 96134 276618
rect 95514 240618 95546 241174
rect 96102 240618 96134 241174
rect 95514 205174 96134 240618
rect 95514 204618 95546 205174
rect 96102 204618 96134 205174
rect 95514 169174 96134 204618
rect 95514 168618 95546 169174
rect 96102 168618 96134 169174
rect 95514 133174 96134 168618
rect 95514 132618 95546 133174
rect 96102 132618 96134 133174
rect 95514 97174 96134 132618
rect 95514 96618 95546 97174
rect 96102 96618 96134 97174
rect 95514 61174 96134 96618
rect 95514 60618 95546 61174
rect 96102 60618 96134 61174
rect 95514 25174 96134 60618
rect 95514 24618 95546 25174
rect 96102 24618 96134 25174
rect 95514 -3226 96134 24618
rect 95514 -3782 95546 -3226
rect 96102 -3782 96134 -3226
rect 95514 -3814 96134 -3782
rect 99234 676894 99854 709082
rect 99234 676338 99266 676894
rect 99822 676338 99854 676894
rect 99234 640894 99854 676338
rect 99234 640338 99266 640894
rect 99822 640338 99854 640894
rect 99234 604894 99854 640338
rect 99234 604338 99266 604894
rect 99822 604338 99854 604894
rect 99234 568894 99854 604338
rect 99234 568338 99266 568894
rect 99822 568338 99854 568894
rect 99234 532894 99854 568338
rect 99234 532338 99266 532894
rect 99822 532338 99854 532894
rect 99234 496894 99854 532338
rect 99234 496338 99266 496894
rect 99822 496338 99854 496894
rect 99234 460894 99854 496338
rect 99234 460338 99266 460894
rect 99822 460338 99854 460894
rect 99234 424894 99854 460338
rect 99234 424338 99266 424894
rect 99822 424338 99854 424894
rect 99234 388894 99854 424338
rect 99234 388338 99266 388894
rect 99822 388338 99854 388894
rect 99234 352894 99854 388338
rect 99234 352338 99266 352894
rect 99822 352338 99854 352894
rect 99234 316894 99854 352338
rect 99234 316338 99266 316894
rect 99822 316338 99854 316894
rect 99234 280894 99854 316338
rect 99234 280338 99266 280894
rect 99822 280338 99854 280894
rect 99234 244894 99854 280338
rect 99234 244338 99266 244894
rect 99822 244338 99854 244894
rect 99234 208894 99854 244338
rect 99234 208338 99266 208894
rect 99822 208338 99854 208894
rect 99234 172894 99854 208338
rect 99234 172338 99266 172894
rect 99822 172338 99854 172894
rect 99234 136894 99854 172338
rect 99234 136338 99266 136894
rect 99822 136338 99854 136894
rect 99234 100894 99854 136338
rect 99234 100338 99266 100894
rect 99822 100338 99854 100894
rect 99234 64894 99854 100338
rect 99234 64338 99266 64894
rect 99822 64338 99854 64894
rect 99234 28894 99854 64338
rect 99234 28338 99266 28894
rect 99822 28338 99854 28894
rect 99234 -5146 99854 28338
rect 99234 -5702 99266 -5146
rect 99822 -5702 99854 -5146
rect 99234 -5734 99854 -5702
rect 102954 680614 103574 711002
rect 120954 710598 121574 711590
rect 120954 710042 120986 710598
rect 121542 710042 121574 710598
rect 117234 708678 117854 709670
rect 117234 708122 117266 708678
rect 117822 708122 117854 708678
rect 113514 706758 114134 707750
rect 113514 706202 113546 706758
rect 114102 706202 114134 706758
rect 102954 680058 102986 680614
rect 103542 680058 103574 680614
rect 102954 644614 103574 680058
rect 102954 644058 102986 644614
rect 103542 644058 103574 644614
rect 102954 608614 103574 644058
rect 102954 608058 102986 608614
rect 103542 608058 103574 608614
rect 102954 572614 103574 608058
rect 102954 572058 102986 572614
rect 103542 572058 103574 572614
rect 102954 536614 103574 572058
rect 102954 536058 102986 536614
rect 103542 536058 103574 536614
rect 102954 500614 103574 536058
rect 102954 500058 102986 500614
rect 103542 500058 103574 500614
rect 102954 464614 103574 500058
rect 102954 464058 102986 464614
rect 103542 464058 103574 464614
rect 102954 428614 103574 464058
rect 102954 428058 102986 428614
rect 103542 428058 103574 428614
rect 102954 392614 103574 428058
rect 102954 392058 102986 392614
rect 103542 392058 103574 392614
rect 102954 356614 103574 392058
rect 102954 356058 102986 356614
rect 103542 356058 103574 356614
rect 102954 320614 103574 356058
rect 102954 320058 102986 320614
rect 103542 320058 103574 320614
rect 102954 284614 103574 320058
rect 102954 284058 102986 284614
rect 103542 284058 103574 284614
rect 102954 248614 103574 284058
rect 102954 248058 102986 248614
rect 103542 248058 103574 248614
rect 102954 212614 103574 248058
rect 102954 212058 102986 212614
rect 103542 212058 103574 212614
rect 102954 176614 103574 212058
rect 102954 176058 102986 176614
rect 103542 176058 103574 176614
rect 102954 140614 103574 176058
rect 102954 140058 102986 140614
rect 103542 140058 103574 140614
rect 102954 104614 103574 140058
rect 102954 104058 102986 104614
rect 103542 104058 103574 104614
rect 102954 68614 103574 104058
rect 102954 68058 102986 68614
rect 103542 68058 103574 68614
rect 102954 32614 103574 68058
rect 102954 32058 102986 32614
rect 103542 32058 103574 32614
rect 84954 -6662 84986 -6106
rect 85542 -6662 85574 -6106
rect 84954 -7654 85574 -6662
rect 102954 -7066 103574 32058
rect 109794 704838 110414 705830
rect 109794 704282 109826 704838
rect 110382 704282 110414 704838
rect 109794 687454 110414 704282
rect 109794 686898 109826 687454
rect 110382 686898 110414 687454
rect 109794 651454 110414 686898
rect 109794 650898 109826 651454
rect 110382 650898 110414 651454
rect 109794 615454 110414 650898
rect 109794 614898 109826 615454
rect 110382 614898 110414 615454
rect 109794 579454 110414 614898
rect 109794 578898 109826 579454
rect 110382 578898 110414 579454
rect 109794 543454 110414 578898
rect 109794 542898 109826 543454
rect 110382 542898 110414 543454
rect 109794 507454 110414 542898
rect 109794 506898 109826 507454
rect 110382 506898 110414 507454
rect 109794 471454 110414 506898
rect 109794 470898 109826 471454
rect 110382 470898 110414 471454
rect 109794 435454 110414 470898
rect 109794 434898 109826 435454
rect 110382 434898 110414 435454
rect 109794 399454 110414 434898
rect 109794 398898 109826 399454
rect 110382 398898 110414 399454
rect 109794 363454 110414 398898
rect 109794 362898 109826 363454
rect 110382 362898 110414 363454
rect 109794 327454 110414 362898
rect 109794 326898 109826 327454
rect 110382 326898 110414 327454
rect 109794 291454 110414 326898
rect 109794 290898 109826 291454
rect 110382 290898 110414 291454
rect 109794 255454 110414 290898
rect 109794 254898 109826 255454
rect 110382 254898 110414 255454
rect 109794 219454 110414 254898
rect 109794 218898 109826 219454
rect 110382 218898 110414 219454
rect 109794 183454 110414 218898
rect 109794 182898 109826 183454
rect 110382 182898 110414 183454
rect 109794 147454 110414 182898
rect 109794 146898 109826 147454
rect 110382 146898 110414 147454
rect 109794 111454 110414 146898
rect 109794 110898 109826 111454
rect 110382 110898 110414 111454
rect 109794 75454 110414 110898
rect 109794 74898 109826 75454
rect 110382 74898 110414 75454
rect 109794 39454 110414 74898
rect 109794 38898 109826 39454
rect 110382 38898 110414 39454
rect 109794 3454 110414 38898
rect 109794 2898 109826 3454
rect 110382 2898 110414 3454
rect 109794 -346 110414 2898
rect 109794 -902 109826 -346
rect 110382 -902 110414 -346
rect 109794 -1894 110414 -902
rect 113514 691174 114134 706202
rect 113514 690618 113546 691174
rect 114102 690618 114134 691174
rect 113514 655174 114134 690618
rect 113514 654618 113546 655174
rect 114102 654618 114134 655174
rect 113514 619174 114134 654618
rect 113514 618618 113546 619174
rect 114102 618618 114134 619174
rect 113514 583174 114134 618618
rect 113514 582618 113546 583174
rect 114102 582618 114134 583174
rect 113514 547174 114134 582618
rect 113514 546618 113546 547174
rect 114102 546618 114134 547174
rect 113514 511174 114134 546618
rect 113514 510618 113546 511174
rect 114102 510618 114134 511174
rect 113514 475174 114134 510618
rect 113514 474618 113546 475174
rect 114102 474618 114134 475174
rect 113514 439174 114134 474618
rect 113514 438618 113546 439174
rect 114102 438618 114134 439174
rect 113514 403174 114134 438618
rect 113514 402618 113546 403174
rect 114102 402618 114134 403174
rect 113514 367174 114134 402618
rect 113514 366618 113546 367174
rect 114102 366618 114134 367174
rect 113514 331174 114134 366618
rect 113514 330618 113546 331174
rect 114102 330618 114134 331174
rect 113514 295174 114134 330618
rect 113514 294618 113546 295174
rect 114102 294618 114134 295174
rect 113514 259174 114134 294618
rect 113514 258618 113546 259174
rect 114102 258618 114134 259174
rect 113514 223174 114134 258618
rect 113514 222618 113546 223174
rect 114102 222618 114134 223174
rect 113514 187174 114134 222618
rect 113514 186618 113546 187174
rect 114102 186618 114134 187174
rect 113514 151174 114134 186618
rect 113514 150618 113546 151174
rect 114102 150618 114134 151174
rect 113514 115174 114134 150618
rect 113514 114618 113546 115174
rect 114102 114618 114134 115174
rect 113514 79174 114134 114618
rect 113514 78618 113546 79174
rect 114102 78618 114134 79174
rect 113514 43174 114134 78618
rect 113514 42618 113546 43174
rect 114102 42618 114134 43174
rect 113514 7174 114134 42618
rect 113514 6618 113546 7174
rect 114102 6618 114134 7174
rect 113514 -2266 114134 6618
rect 113514 -2822 113546 -2266
rect 114102 -2822 114134 -2266
rect 113514 -3814 114134 -2822
rect 117234 694894 117854 708122
rect 117234 694338 117266 694894
rect 117822 694338 117854 694894
rect 117234 658894 117854 694338
rect 117234 658338 117266 658894
rect 117822 658338 117854 658894
rect 117234 622894 117854 658338
rect 117234 622338 117266 622894
rect 117822 622338 117854 622894
rect 117234 586894 117854 622338
rect 117234 586338 117266 586894
rect 117822 586338 117854 586894
rect 117234 550894 117854 586338
rect 117234 550338 117266 550894
rect 117822 550338 117854 550894
rect 117234 514894 117854 550338
rect 117234 514338 117266 514894
rect 117822 514338 117854 514894
rect 117234 478894 117854 514338
rect 117234 478338 117266 478894
rect 117822 478338 117854 478894
rect 117234 442894 117854 478338
rect 117234 442338 117266 442894
rect 117822 442338 117854 442894
rect 117234 406894 117854 442338
rect 117234 406338 117266 406894
rect 117822 406338 117854 406894
rect 117234 370894 117854 406338
rect 117234 370338 117266 370894
rect 117822 370338 117854 370894
rect 117234 334894 117854 370338
rect 117234 334338 117266 334894
rect 117822 334338 117854 334894
rect 117234 298894 117854 334338
rect 117234 298338 117266 298894
rect 117822 298338 117854 298894
rect 117234 262894 117854 298338
rect 117234 262338 117266 262894
rect 117822 262338 117854 262894
rect 117234 226894 117854 262338
rect 117234 226338 117266 226894
rect 117822 226338 117854 226894
rect 117234 190894 117854 226338
rect 117234 190338 117266 190894
rect 117822 190338 117854 190894
rect 117234 154894 117854 190338
rect 117234 154338 117266 154894
rect 117822 154338 117854 154894
rect 117234 118894 117854 154338
rect 117234 118338 117266 118894
rect 117822 118338 117854 118894
rect 117234 82894 117854 118338
rect 117234 82338 117266 82894
rect 117822 82338 117854 82894
rect 117234 46894 117854 82338
rect 117234 46338 117266 46894
rect 117822 46338 117854 46894
rect 117234 10894 117854 46338
rect 117234 10338 117266 10894
rect 117822 10338 117854 10894
rect 117234 -4186 117854 10338
rect 117234 -4742 117266 -4186
rect 117822 -4742 117854 -4186
rect 117234 -5734 117854 -4742
rect 120954 698614 121574 710042
rect 138954 711558 139574 711590
rect 138954 711002 138986 711558
rect 139542 711002 139574 711558
rect 135234 709638 135854 709670
rect 135234 709082 135266 709638
rect 135822 709082 135854 709638
rect 131514 707718 132134 707750
rect 131514 707162 131546 707718
rect 132102 707162 132134 707718
rect 120954 698058 120986 698614
rect 121542 698058 121574 698614
rect 120954 662614 121574 698058
rect 120954 662058 120986 662614
rect 121542 662058 121574 662614
rect 120954 626614 121574 662058
rect 120954 626058 120986 626614
rect 121542 626058 121574 626614
rect 120954 590614 121574 626058
rect 120954 590058 120986 590614
rect 121542 590058 121574 590614
rect 120954 554614 121574 590058
rect 120954 554058 120986 554614
rect 121542 554058 121574 554614
rect 120954 518614 121574 554058
rect 120954 518058 120986 518614
rect 121542 518058 121574 518614
rect 120954 482614 121574 518058
rect 120954 482058 120986 482614
rect 121542 482058 121574 482614
rect 120954 446614 121574 482058
rect 120954 446058 120986 446614
rect 121542 446058 121574 446614
rect 120954 410614 121574 446058
rect 120954 410058 120986 410614
rect 121542 410058 121574 410614
rect 120954 374614 121574 410058
rect 120954 374058 120986 374614
rect 121542 374058 121574 374614
rect 120954 338614 121574 374058
rect 120954 338058 120986 338614
rect 121542 338058 121574 338614
rect 120954 302614 121574 338058
rect 120954 302058 120986 302614
rect 121542 302058 121574 302614
rect 120954 266614 121574 302058
rect 120954 266058 120986 266614
rect 121542 266058 121574 266614
rect 120954 230614 121574 266058
rect 120954 230058 120986 230614
rect 121542 230058 121574 230614
rect 120954 194614 121574 230058
rect 120954 194058 120986 194614
rect 121542 194058 121574 194614
rect 120954 158614 121574 194058
rect 120954 158058 120986 158614
rect 121542 158058 121574 158614
rect 120954 122614 121574 158058
rect 120954 122058 120986 122614
rect 121542 122058 121574 122614
rect 120954 86614 121574 122058
rect 120954 86058 120986 86614
rect 121542 86058 121574 86614
rect 120954 50614 121574 86058
rect 120954 50058 120986 50614
rect 121542 50058 121574 50614
rect 120954 14614 121574 50058
rect 120954 14058 120986 14614
rect 121542 14058 121574 14614
rect 102954 -7622 102986 -7066
rect 103542 -7622 103574 -7066
rect 102954 -7654 103574 -7622
rect 120954 -6106 121574 14058
rect 127794 705798 128414 705830
rect 127794 705242 127826 705798
rect 128382 705242 128414 705798
rect 127794 669454 128414 705242
rect 127794 668898 127826 669454
rect 128382 668898 128414 669454
rect 127794 633454 128414 668898
rect 127794 632898 127826 633454
rect 128382 632898 128414 633454
rect 127794 597454 128414 632898
rect 127794 596898 127826 597454
rect 128382 596898 128414 597454
rect 127794 561454 128414 596898
rect 127794 560898 127826 561454
rect 128382 560898 128414 561454
rect 127794 525454 128414 560898
rect 127794 524898 127826 525454
rect 128382 524898 128414 525454
rect 127794 489454 128414 524898
rect 127794 488898 127826 489454
rect 128382 488898 128414 489454
rect 127794 453454 128414 488898
rect 127794 452898 127826 453454
rect 128382 452898 128414 453454
rect 127794 417454 128414 452898
rect 127794 416898 127826 417454
rect 128382 416898 128414 417454
rect 127794 381454 128414 416898
rect 127794 380898 127826 381454
rect 128382 380898 128414 381454
rect 127794 345454 128414 380898
rect 127794 344898 127826 345454
rect 128382 344898 128414 345454
rect 127794 309454 128414 344898
rect 127794 308898 127826 309454
rect 128382 308898 128414 309454
rect 127794 273454 128414 308898
rect 127794 272898 127826 273454
rect 128382 272898 128414 273454
rect 127794 237454 128414 272898
rect 127794 236898 127826 237454
rect 128382 236898 128414 237454
rect 127794 201454 128414 236898
rect 127794 200898 127826 201454
rect 128382 200898 128414 201454
rect 127794 165454 128414 200898
rect 127794 164898 127826 165454
rect 128382 164898 128414 165454
rect 127794 129454 128414 164898
rect 127794 128898 127826 129454
rect 128382 128898 128414 129454
rect 127794 93454 128414 128898
rect 127794 92898 127826 93454
rect 128382 92898 128414 93454
rect 127794 57454 128414 92898
rect 127794 56898 127826 57454
rect 128382 56898 128414 57454
rect 127794 21454 128414 56898
rect 127794 20898 127826 21454
rect 128382 20898 128414 21454
rect 127794 -1306 128414 20898
rect 127794 -1862 127826 -1306
rect 128382 -1862 128414 -1306
rect 127794 -1894 128414 -1862
rect 131514 673174 132134 707162
rect 131514 672618 131546 673174
rect 132102 672618 132134 673174
rect 131514 637174 132134 672618
rect 131514 636618 131546 637174
rect 132102 636618 132134 637174
rect 131514 601174 132134 636618
rect 131514 600618 131546 601174
rect 132102 600618 132134 601174
rect 131514 565174 132134 600618
rect 131514 564618 131546 565174
rect 132102 564618 132134 565174
rect 131514 529174 132134 564618
rect 131514 528618 131546 529174
rect 132102 528618 132134 529174
rect 131514 493174 132134 528618
rect 131514 492618 131546 493174
rect 132102 492618 132134 493174
rect 131514 457174 132134 492618
rect 131514 456618 131546 457174
rect 132102 456618 132134 457174
rect 131514 421174 132134 456618
rect 131514 420618 131546 421174
rect 132102 420618 132134 421174
rect 131514 385174 132134 420618
rect 131514 384618 131546 385174
rect 132102 384618 132134 385174
rect 131514 349174 132134 384618
rect 131514 348618 131546 349174
rect 132102 348618 132134 349174
rect 131514 313174 132134 348618
rect 131514 312618 131546 313174
rect 132102 312618 132134 313174
rect 131514 277174 132134 312618
rect 131514 276618 131546 277174
rect 132102 276618 132134 277174
rect 131514 241174 132134 276618
rect 131514 240618 131546 241174
rect 132102 240618 132134 241174
rect 131514 205174 132134 240618
rect 131514 204618 131546 205174
rect 132102 204618 132134 205174
rect 131514 169174 132134 204618
rect 131514 168618 131546 169174
rect 132102 168618 132134 169174
rect 131514 133174 132134 168618
rect 131514 132618 131546 133174
rect 132102 132618 132134 133174
rect 131514 97174 132134 132618
rect 131514 96618 131546 97174
rect 132102 96618 132134 97174
rect 131514 61174 132134 96618
rect 131514 60618 131546 61174
rect 132102 60618 132134 61174
rect 131514 25174 132134 60618
rect 131514 24618 131546 25174
rect 132102 24618 132134 25174
rect 131514 -3226 132134 24618
rect 131514 -3782 131546 -3226
rect 132102 -3782 132134 -3226
rect 131514 -3814 132134 -3782
rect 135234 676894 135854 709082
rect 135234 676338 135266 676894
rect 135822 676338 135854 676894
rect 135234 640894 135854 676338
rect 135234 640338 135266 640894
rect 135822 640338 135854 640894
rect 135234 604894 135854 640338
rect 135234 604338 135266 604894
rect 135822 604338 135854 604894
rect 135234 568894 135854 604338
rect 135234 568338 135266 568894
rect 135822 568338 135854 568894
rect 135234 532894 135854 568338
rect 135234 532338 135266 532894
rect 135822 532338 135854 532894
rect 135234 496894 135854 532338
rect 135234 496338 135266 496894
rect 135822 496338 135854 496894
rect 135234 460894 135854 496338
rect 135234 460338 135266 460894
rect 135822 460338 135854 460894
rect 135234 424894 135854 460338
rect 135234 424338 135266 424894
rect 135822 424338 135854 424894
rect 135234 388894 135854 424338
rect 135234 388338 135266 388894
rect 135822 388338 135854 388894
rect 135234 352894 135854 388338
rect 135234 352338 135266 352894
rect 135822 352338 135854 352894
rect 135234 316894 135854 352338
rect 135234 316338 135266 316894
rect 135822 316338 135854 316894
rect 135234 280894 135854 316338
rect 135234 280338 135266 280894
rect 135822 280338 135854 280894
rect 135234 244894 135854 280338
rect 135234 244338 135266 244894
rect 135822 244338 135854 244894
rect 135234 208894 135854 244338
rect 135234 208338 135266 208894
rect 135822 208338 135854 208894
rect 135234 172894 135854 208338
rect 135234 172338 135266 172894
rect 135822 172338 135854 172894
rect 135234 136894 135854 172338
rect 135234 136338 135266 136894
rect 135822 136338 135854 136894
rect 135234 100894 135854 136338
rect 135234 100338 135266 100894
rect 135822 100338 135854 100894
rect 135234 64894 135854 100338
rect 135234 64338 135266 64894
rect 135822 64338 135854 64894
rect 135234 28894 135854 64338
rect 135234 28338 135266 28894
rect 135822 28338 135854 28894
rect 135234 -5146 135854 28338
rect 135234 -5702 135266 -5146
rect 135822 -5702 135854 -5146
rect 135234 -5734 135854 -5702
rect 138954 680614 139574 711002
rect 156954 710598 157574 711590
rect 156954 710042 156986 710598
rect 157542 710042 157574 710598
rect 153234 708678 153854 709670
rect 153234 708122 153266 708678
rect 153822 708122 153854 708678
rect 149514 706758 150134 707750
rect 149514 706202 149546 706758
rect 150102 706202 150134 706758
rect 138954 680058 138986 680614
rect 139542 680058 139574 680614
rect 138954 644614 139574 680058
rect 138954 644058 138986 644614
rect 139542 644058 139574 644614
rect 138954 608614 139574 644058
rect 138954 608058 138986 608614
rect 139542 608058 139574 608614
rect 138954 572614 139574 608058
rect 138954 572058 138986 572614
rect 139542 572058 139574 572614
rect 138954 536614 139574 572058
rect 138954 536058 138986 536614
rect 139542 536058 139574 536614
rect 138954 500614 139574 536058
rect 138954 500058 138986 500614
rect 139542 500058 139574 500614
rect 138954 464614 139574 500058
rect 138954 464058 138986 464614
rect 139542 464058 139574 464614
rect 138954 428614 139574 464058
rect 138954 428058 138986 428614
rect 139542 428058 139574 428614
rect 138954 392614 139574 428058
rect 138954 392058 138986 392614
rect 139542 392058 139574 392614
rect 138954 356614 139574 392058
rect 138954 356058 138986 356614
rect 139542 356058 139574 356614
rect 138954 320614 139574 356058
rect 138954 320058 138986 320614
rect 139542 320058 139574 320614
rect 138954 284614 139574 320058
rect 138954 284058 138986 284614
rect 139542 284058 139574 284614
rect 138954 248614 139574 284058
rect 138954 248058 138986 248614
rect 139542 248058 139574 248614
rect 138954 212614 139574 248058
rect 138954 212058 138986 212614
rect 139542 212058 139574 212614
rect 138954 176614 139574 212058
rect 138954 176058 138986 176614
rect 139542 176058 139574 176614
rect 138954 140614 139574 176058
rect 138954 140058 138986 140614
rect 139542 140058 139574 140614
rect 138954 104614 139574 140058
rect 138954 104058 138986 104614
rect 139542 104058 139574 104614
rect 138954 68614 139574 104058
rect 138954 68058 138986 68614
rect 139542 68058 139574 68614
rect 138954 32614 139574 68058
rect 138954 32058 138986 32614
rect 139542 32058 139574 32614
rect 120954 -6662 120986 -6106
rect 121542 -6662 121574 -6106
rect 120954 -7654 121574 -6662
rect 138954 -7066 139574 32058
rect 145794 704838 146414 705830
rect 145794 704282 145826 704838
rect 146382 704282 146414 704838
rect 145794 687454 146414 704282
rect 145794 686898 145826 687454
rect 146382 686898 146414 687454
rect 145794 651454 146414 686898
rect 145794 650898 145826 651454
rect 146382 650898 146414 651454
rect 145794 615454 146414 650898
rect 145794 614898 145826 615454
rect 146382 614898 146414 615454
rect 145794 579454 146414 614898
rect 145794 578898 145826 579454
rect 146382 578898 146414 579454
rect 145794 543454 146414 578898
rect 145794 542898 145826 543454
rect 146382 542898 146414 543454
rect 145794 507454 146414 542898
rect 145794 506898 145826 507454
rect 146382 506898 146414 507454
rect 145794 471454 146414 506898
rect 145794 470898 145826 471454
rect 146382 470898 146414 471454
rect 145794 435454 146414 470898
rect 145794 434898 145826 435454
rect 146382 434898 146414 435454
rect 145794 399454 146414 434898
rect 145794 398898 145826 399454
rect 146382 398898 146414 399454
rect 145794 363454 146414 398898
rect 145794 362898 145826 363454
rect 146382 362898 146414 363454
rect 145794 327454 146414 362898
rect 145794 326898 145826 327454
rect 146382 326898 146414 327454
rect 145794 291454 146414 326898
rect 145794 290898 145826 291454
rect 146382 290898 146414 291454
rect 145794 255454 146414 290898
rect 145794 254898 145826 255454
rect 146382 254898 146414 255454
rect 145794 219454 146414 254898
rect 145794 218898 145826 219454
rect 146382 218898 146414 219454
rect 145794 183454 146414 218898
rect 145794 182898 145826 183454
rect 146382 182898 146414 183454
rect 145794 147454 146414 182898
rect 145794 146898 145826 147454
rect 146382 146898 146414 147454
rect 145794 111454 146414 146898
rect 145794 110898 145826 111454
rect 146382 110898 146414 111454
rect 145794 75454 146414 110898
rect 145794 74898 145826 75454
rect 146382 74898 146414 75454
rect 145794 39454 146414 74898
rect 145794 38898 145826 39454
rect 146382 38898 146414 39454
rect 145794 3454 146414 38898
rect 145794 2898 145826 3454
rect 146382 2898 146414 3454
rect 145794 -346 146414 2898
rect 145794 -902 145826 -346
rect 146382 -902 146414 -346
rect 145794 -1894 146414 -902
rect 149514 691174 150134 706202
rect 149514 690618 149546 691174
rect 150102 690618 150134 691174
rect 149514 655174 150134 690618
rect 149514 654618 149546 655174
rect 150102 654618 150134 655174
rect 149514 619174 150134 654618
rect 149514 618618 149546 619174
rect 150102 618618 150134 619174
rect 149514 583174 150134 618618
rect 149514 582618 149546 583174
rect 150102 582618 150134 583174
rect 149514 547174 150134 582618
rect 149514 546618 149546 547174
rect 150102 546618 150134 547174
rect 149514 511174 150134 546618
rect 149514 510618 149546 511174
rect 150102 510618 150134 511174
rect 149514 475174 150134 510618
rect 149514 474618 149546 475174
rect 150102 474618 150134 475174
rect 149514 439174 150134 474618
rect 149514 438618 149546 439174
rect 150102 438618 150134 439174
rect 149514 403174 150134 438618
rect 149514 402618 149546 403174
rect 150102 402618 150134 403174
rect 149514 367174 150134 402618
rect 149514 366618 149546 367174
rect 150102 366618 150134 367174
rect 149514 331174 150134 366618
rect 149514 330618 149546 331174
rect 150102 330618 150134 331174
rect 149514 295174 150134 330618
rect 149514 294618 149546 295174
rect 150102 294618 150134 295174
rect 149514 259174 150134 294618
rect 149514 258618 149546 259174
rect 150102 258618 150134 259174
rect 149514 223174 150134 258618
rect 149514 222618 149546 223174
rect 150102 222618 150134 223174
rect 149514 187174 150134 222618
rect 149514 186618 149546 187174
rect 150102 186618 150134 187174
rect 149514 151174 150134 186618
rect 149514 150618 149546 151174
rect 150102 150618 150134 151174
rect 149514 115174 150134 150618
rect 149514 114618 149546 115174
rect 150102 114618 150134 115174
rect 149514 79174 150134 114618
rect 149514 78618 149546 79174
rect 150102 78618 150134 79174
rect 149514 43174 150134 78618
rect 149514 42618 149546 43174
rect 150102 42618 150134 43174
rect 149514 7174 150134 42618
rect 149514 6618 149546 7174
rect 150102 6618 150134 7174
rect 149514 -2266 150134 6618
rect 149514 -2822 149546 -2266
rect 150102 -2822 150134 -2266
rect 149514 -3814 150134 -2822
rect 153234 694894 153854 708122
rect 153234 694338 153266 694894
rect 153822 694338 153854 694894
rect 153234 658894 153854 694338
rect 153234 658338 153266 658894
rect 153822 658338 153854 658894
rect 153234 622894 153854 658338
rect 153234 622338 153266 622894
rect 153822 622338 153854 622894
rect 153234 586894 153854 622338
rect 153234 586338 153266 586894
rect 153822 586338 153854 586894
rect 153234 550894 153854 586338
rect 153234 550338 153266 550894
rect 153822 550338 153854 550894
rect 153234 514894 153854 550338
rect 153234 514338 153266 514894
rect 153822 514338 153854 514894
rect 153234 478894 153854 514338
rect 153234 478338 153266 478894
rect 153822 478338 153854 478894
rect 153234 442894 153854 478338
rect 153234 442338 153266 442894
rect 153822 442338 153854 442894
rect 153234 406894 153854 442338
rect 153234 406338 153266 406894
rect 153822 406338 153854 406894
rect 153234 370894 153854 406338
rect 153234 370338 153266 370894
rect 153822 370338 153854 370894
rect 153234 334894 153854 370338
rect 153234 334338 153266 334894
rect 153822 334338 153854 334894
rect 153234 298894 153854 334338
rect 153234 298338 153266 298894
rect 153822 298338 153854 298894
rect 153234 262894 153854 298338
rect 153234 262338 153266 262894
rect 153822 262338 153854 262894
rect 153234 226894 153854 262338
rect 153234 226338 153266 226894
rect 153822 226338 153854 226894
rect 153234 190894 153854 226338
rect 153234 190338 153266 190894
rect 153822 190338 153854 190894
rect 153234 154894 153854 190338
rect 153234 154338 153266 154894
rect 153822 154338 153854 154894
rect 153234 118894 153854 154338
rect 153234 118338 153266 118894
rect 153822 118338 153854 118894
rect 153234 82894 153854 118338
rect 153234 82338 153266 82894
rect 153822 82338 153854 82894
rect 153234 46894 153854 82338
rect 153234 46338 153266 46894
rect 153822 46338 153854 46894
rect 153234 10894 153854 46338
rect 153234 10338 153266 10894
rect 153822 10338 153854 10894
rect 153234 -4186 153854 10338
rect 153234 -4742 153266 -4186
rect 153822 -4742 153854 -4186
rect 153234 -5734 153854 -4742
rect 156954 698614 157574 710042
rect 174954 711558 175574 711590
rect 174954 711002 174986 711558
rect 175542 711002 175574 711558
rect 171234 709638 171854 709670
rect 171234 709082 171266 709638
rect 171822 709082 171854 709638
rect 167514 707718 168134 707750
rect 167514 707162 167546 707718
rect 168102 707162 168134 707718
rect 156954 698058 156986 698614
rect 157542 698058 157574 698614
rect 156954 662614 157574 698058
rect 156954 662058 156986 662614
rect 157542 662058 157574 662614
rect 156954 626614 157574 662058
rect 156954 626058 156986 626614
rect 157542 626058 157574 626614
rect 156954 590614 157574 626058
rect 156954 590058 156986 590614
rect 157542 590058 157574 590614
rect 156954 554614 157574 590058
rect 156954 554058 156986 554614
rect 157542 554058 157574 554614
rect 156954 518614 157574 554058
rect 156954 518058 156986 518614
rect 157542 518058 157574 518614
rect 156954 482614 157574 518058
rect 156954 482058 156986 482614
rect 157542 482058 157574 482614
rect 156954 446614 157574 482058
rect 156954 446058 156986 446614
rect 157542 446058 157574 446614
rect 156954 410614 157574 446058
rect 156954 410058 156986 410614
rect 157542 410058 157574 410614
rect 156954 374614 157574 410058
rect 156954 374058 156986 374614
rect 157542 374058 157574 374614
rect 156954 338614 157574 374058
rect 156954 338058 156986 338614
rect 157542 338058 157574 338614
rect 156954 302614 157574 338058
rect 156954 302058 156986 302614
rect 157542 302058 157574 302614
rect 156954 266614 157574 302058
rect 156954 266058 156986 266614
rect 157542 266058 157574 266614
rect 156954 230614 157574 266058
rect 156954 230058 156986 230614
rect 157542 230058 157574 230614
rect 156954 194614 157574 230058
rect 156954 194058 156986 194614
rect 157542 194058 157574 194614
rect 156954 158614 157574 194058
rect 156954 158058 156986 158614
rect 157542 158058 157574 158614
rect 156954 122614 157574 158058
rect 156954 122058 156986 122614
rect 157542 122058 157574 122614
rect 156954 86614 157574 122058
rect 156954 86058 156986 86614
rect 157542 86058 157574 86614
rect 156954 50614 157574 86058
rect 156954 50058 156986 50614
rect 157542 50058 157574 50614
rect 156954 14614 157574 50058
rect 156954 14058 156986 14614
rect 157542 14058 157574 14614
rect 138954 -7622 138986 -7066
rect 139542 -7622 139574 -7066
rect 138954 -7654 139574 -7622
rect 156954 -6106 157574 14058
rect 163794 705798 164414 705830
rect 163794 705242 163826 705798
rect 164382 705242 164414 705798
rect 163794 669454 164414 705242
rect 163794 668898 163826 669454
rect 164382 668898 164414 669454
rect 163794 633454 164414 668898
rect 163794 632898 163826 633454
rect 164382 632898 164414 633454
rect 163794 597454 164414 632898
rect 163794 596898 163826 597454
rect 164382 596898 164414 597454
rect 163794 561454 164414 596898
rect 163794 560898 163826 561454
rect 164382 560898 164414 561454
rect 163794 525454 164414 560898
rect 163794 524898 163826 525454
rect 164382 524898 164414 525454
rect 163794 489454 164414 524898
rect 163794 488898 163826 489454
rect 164382 488898 164414 489454
rect 163794 453454 164414 488898
rect 163794 452898 163826 453454
rect 164382 452898 164414 453454
rect 163794 417454 164414 452898
rect 163794 416898 163826 417454
rect 164382 416898 164414 417454
rect 163794 381454 164414 416898
rect 163794 380898 163826 381454
rect 164382 380898 164414 381454
rect 163794 345454 164414 380898
rect 163794 344898 163826 345454
rect 164382 344898 164414 345454
rect 163794 309454 164414 344898
rect 163794 308898 163826 309454
rect 164382 308898 164414 309454
rect 163794 273454 164414 308898
rect 163794 272898 163826 273454
rect 164382 272898 164414 273454
rect 163794 237454 164414 272898
rect 163794 236898 163826 237454
rect 164382 236898 164414 237454
rect 163794 201454 164414 236898
rect 163794 200898 163826 201454
rect 164382 200898 164414 201454
rect 163794 165454 164414 200898
rect 163794 164898 163826 165454
rect 164382 164898 164414 165454
rect 163794 129454 164414 164898
rect 163794 128898 163826 129454
rect 164382 128898 164414 129454
rect 163794 93454 164414 128898
rect 163794 92898 163826 93454
rect 164382 92898 164414 93454
rect 163794 57454 164414 92898
rect 163794 56898 163826 57454
rect 164382 56898 164414 57454
rect 163794 21454 164414 56898
rect 163794 20898 163826 21454
rect 164382 20898 164414 21454
rect 163794 -1306 164414 20898
rect 163794 -1862 163826 -1306
rect 164382 -1862 164414 -1306
rect 163794 -1894 164414 -1862
rect 167514 673174 168134 707162
rect 167514 672618 167546 673174
rect 168102 672618 168134 673174
rect 167514 637174 168134 672618
rect 167514 636618 167546 637174
rect 168102 636618 168134 637174
rect 167514 601174 168134 636618
rect 167514 600618 167546 601174
rect 168102 600618 168134 601174
rect 167514 565174 168134 600618
rect 167514 564618 167546 565174
rect 168102 564618 168134 565174
rect 167514 529174 168134 564618
rect 167514 528618 167546 529174
rect 168102 528618 168134 529174
rect 167514 493174 168134 528618
rect 167514 492618 167546 493174
rect 168102 492618 168134 493174
rect 167514 457174 168134 492618
rect 167514 456618 167546 457174
rect 168102 456618 168134 457174
rect 167514 421174 168134 456618
rect 167514 420618 167546 421174
rect 168102 420618 168134 421174
rect 167514 385174 168134 420618
rect 167514 384618 167546 385174
rect 168102 384618 168134 385174
rect 167514 349174 168134 384618
rect 167514 348618 167546 349174
rect 168102 348618 168134 349174
rect 167514 313174 168134 348618
rect 167514 312618 167546 313174
rect 168102 312618 168134 313174
rect 167514 277174 168134 312618
rect 167514 276618 167546 277174
rect 168102 276618 168134 277174
rect 167514 241174 168134 276618
rect 167514 240618 167546 241174
rect 168102 240618 168134 241174
rect 167514 205174 168134 240618
rect 167514 204618 167546 205174
rect 168102 204618 168134 205174
rect 167514 169174 168134 204618
rect 167514 168618 167546 169174
rect 168102 168618 168134 169174
rect 167514 133174 168134 168618
rect 167514 132618 167546 133174
rect 168102 132618 168134 133174
rect 167514 97174 168134 132618
rect 167514 96618 167546 97174
rect 168102 96618 168134 97174
rect 167514 61174 168134 96618
rect 167514 60618 167546 61174
rect 168102 60618 168134 61174
rect 167514 25174 168134 60618
rect 167514 24618 167546 25174
rect 168102 24618 168134 25174
rect 167514 -3226 168134 24618
rect 167514 -3782 167546 -3226
rect 168102 -3782 168134 -3226
rect 167514 -3814 168134 -3782
rect 171234 676894 171854 709082
rect 171234 676338 171266 676894
rect 171822 676338 171854 676894
rect 171234 640894 171854 676338
rect 171234 640338 171266 640894
rect 171822 640338 171854 640894
rect 171234 604894 171854 640338
rect 171234 604338 171266 604894
rect 171822 604338 171854 604894
rect 171234 568894 171854 604338
rect 171234 568338 171266 568894
rect 171822 568338 171854 568894
rect 171234 532894 171854 568338
rect 171234 532338 171266 532894
rect 171822 532338 171854 532894
rect 171234 496894 171854 532338
rect 171234 496338 171266 496894
rect 171822 496338 171854 496894
rect 171234 460894 171854 496338
rect 171234 460338 171266 460894
rect 171822 460338 171854 460894
rect 171234 424894 171854 460338
rect 171234 424338 171266 424894
rect 171822 424338 171854 424894
rect 171234 388894 171854 424338
rect 171234 388338 171266 388894
rect 171822 388338 171854 388894
rect 171234 352894 171854 388338
rect 171234 352338 171266 352894
rect 171822 352338 171854 352894
rect 171234 316894 171854 352338
rect 171234 316338 171266 316894
rect 171822 316338 171854 316894
rect 171234 280894 171854 316338
rect 171234 280338 171266 280894
rect 171822 280338 171854 280894
rect 171234 244894 171854 280338
rect 171234 244338 171266 244894
rect 171822 244338 171854 244894
rect 171234 208894 171854 244338
rect 171234 208338 171266 208894
rect 171822 208338 171854 208894
rect 171234 172894 171854 208338
rect 171234 172338 171266 172894
rect 171822 172338 171854 172894
rect 171234 136894 171854 172338
rect 171234 136338 171266 136894
rect 171822 136338 171854 136894
rect 171234 100894 171854 136338
rect 171234 100338 171266 100894
rect 171822 100338 171854 100894
rect 171234 64894 171854 100338
rect 171234 64338 171266 64894
rect 171822 64338 171854 64894
rect 171234 28894 171854 64338
rect 171234 28338 171266 28894
rect 171822 28338 171854 28894
rect 171234 -5146 171854 28338
rect 171234 -5702 171266 -5146
rect 171822 -5702 171854 -5146
rect 171234 -5734 171854 -5702
rect 174954 680614 175574 711002
rect 192954 710598 193574 711590
rect 192954 710042 192986 710598
rect 193542 710042 193574 710598
rect 189234 708678 189854 709670
rect 189234 708122 189266 708678
rect 189822 708122 189854 708678
rect 185514 706758 186134 707750
rect 185514 706202 185546 706758
rect 186102 706202 186134 706758
rect 174954 680058 174986 680614
rect 175542 680058 175574 680614
rect 174954 644614 175574 680058
rect 174954 644058 174986 644614
rect 175542 644058 175574 644614
rect 174954 608614 175574 644058
rect 174954 608058 174986 608614
rect 175542 608058 175574 608614
rect 174954 572614 175574 608058
rect 174954 572058 174986 572614
rect 175542 572058 175574 572614
rect 174954 536614 175574 572058
rect 174954 536058 174986 536614
rect 175542 536058 175574 536614
rect 174954 500614 175574 536058
rect 174954 500058 174986 500614
rect 175542 500058 175574 500614
rect 174954 464614 175574 500058
rect 174954 464058 174986 464614
rect 175542 464058 175574 464614
rect 174954 428614 175574 464058
rect 174954 428058 174986 428614
rect 175542 428058 175574 428614
rect 174954 392614 175574 428058
rect 174954 392058 174986 392614
rect 175542 392058 175574 392614
rect 174954 356614 175574 392058
rect 174954 356058 174986 356614
rect 175542 356058 175574 356614
rect 174954 320614 175574 356058
rect 174954 320058 174986 320614
rect 175542 320058 175574 320614
rect 174954 284614 175574 320058
rect 174954 284058 174986 284614
rect 175542 284058 175574 284614
rect 174954 248614 175574 284058
rect 174954 248058 174986 248614
rect 175542 248058 175574 248614
rect 174954 212614 175574 248058
rect 174954 212058 174986 212614
rect 175542 212058 175574 212614
rect 174954 176614 175574 212058
rect 174954 176058 174986 176614
rect 175542 176058 175574 176614
rect 174954 140614 175574 176058
rect 174954 140058 174986 140614
rect 175542 140058 175574 140614
rect 174954 104614 175574 140058
rect 174954 104058 174986 104614
rect 175542 104058 175574 104614
rect 174954 68614 175574 104058
rect 174954 68058 174986 68614
rect 175542 68058 175574 68614
rect 174954 32614 175574 68058
rect 174954 32058 174986 32614
rect 175542 32058 175574 32614
rect 156954 -6662 156986 -6106
rect 157542 -6662 157574 -6106
rect 156954 -7654 157574 -6662
rect 174954 -7066 175574 32058
rect 181794 704838 182414 705830
rect 181794 704282 181826 704838
rect 182382 704282 182414 704838
rect 181794 687454 182414 704282
rect 181794 686898 181826 687454
rect 182382 686898 182414 687454
rect 181794 651454 182414 686898
rect 181794 650898 181826 651454
rect 182382 650898 182414 651454
rect 181794 615454 182414 650898
rect 181794 614898 181826 615454
rect 182382 614898 182414 615454
rect 181794 579454 182414 614898
rect 181794 578898 181826 579454
rect 182382 578898 182414 579454
rect 181794 543454 182414 578898
rect 181794 542898 181826 543454
rect 182382 542898 182414 543454
rect 181794 507454 182414 542898
rect 181794 506898 181826 507454
rect 182382 506898 182414 507454
rect 181794 471454 182414 506898
rect 181794 470898 181826 471454
rect 182382 470898 182414 471454
rect 181794 435454 182414 470898
rect 181794 434898 181826 435454
rect 182382 434898 182414 435454
rect 181794 399454 182414 434898
rect 181794 398898 181826 399454
rect 182382 398898 182414 399454
rect 181794 363454 182414 398898
rect 181794 362898 181826 363454
rect 182382 362898 182414 363454
rect 181794 327454 182414 362898
rect 181794 326898 181826 327454
rect 182382 326898 182414 327454
rect 181794 291454 182414 326898
rect 181794 290898 181826 291454
rect 182382 290898 182414 291454
rect 181794 255454 182414 290898
rect 181794 254898 181826 255454
rect 182382 254898 182414 255454
rect 181794 219454 182414 254898
rect 181794 218898 181826 219454
rect 182382 218898 182414 219454
rect 181794 183454 182414 218898
rect 181794 182898 181826 183454
rect 182382 182898 182414 183454
rect 181794 147454 182414 182898
rect 181794 146898 181826 147454
rect 182382 146898 182414 147454
rect 181794 111454 182414 146898
rect 181794 110898 181826 111454
rect 182382 110898 182414 111454
rect 181794 75454 182414 110898
rect 181794 74898 181826 75454
rect 182382 74898 182414 75454
rect 181794 39454 182414 74898
rect 181794 38898 181826 39454
rect 182382 38898 182414 39454
rect 181794 3454 182414 38898
rect 181794 2898 181826 3454
rect 182382 2898 182414 3454
rect 181794 -346 182414 2898
rect 181794 -902 181826 -346
rect 182382 -902 182414 -346
rect 181794 -1894 182414 -902
rect 185514 691174 186134 706202
rect 185514 690618 185546 691174
rect 186102 690618 186134 691174
rect 185514 655174 186134 690618
rect 185514 654618 185546 655174
rect 186102 654618 186134 655174
rect 185514 619174 186134 654618
rect 185514 618618 185546 619174
rect 186102 618618 186134 619174
rect 185514 583174 186134 618618
rect 185514 582618 185546 583174
rect 186102 582618 186134 583174
rect 185514 547174 186134 582618
rect 185514 546618 185546 547174
rect 186102 546618 186134 547174
rect 185514 511174 186134 546618
rect 185514 510618 185546 511174
rect 186102 510618 186134 511174
rect 185514 475174 186134 510618
rect 185514 474618 185546 475174
rect 186102 474618 186134 475174
rect 185514 439174 186134 474618
rect 185514 438618 185546 439174
rect 186102 438618 186134 439174
rect 185514 403174 186134 438618
rect 185514 402618 185546 403174
rect 186102 402618 186134 403174
rect 185514 367174 186134 402618
rect 185514 366618 185546 367174
rect 186102 366618 186134 367174
rect 185514 331174 186134 366618
rect 185514 330618 185546 331174
rect 186102 330618 186134 331174
rect 185514 295174 186134 330618
rect 185514 294618 185546 295174
rect 186102 294618 186134 295174
rect 185514 259174 186134 294618
rect 185514 258618 185546 259174
rect 186102 258618 186134 259174
rect 185514 223174 186134 258618
rect 185514 222618 185546 223174
rect 186102 222618 186134 223174
rect 185514 187174 186134 222618
rect 185514 186618 185546 187174
rect 186102 186618 186134 187174
rect 185514 151174 186134 186618
rect 185514 150618 185546 151174
rect 186102 150618 186134 151174
rect 185514 115174 186134 150618
rect 185514 114618 185546 115174
rect 186102 114618 186134 115174
rect 185514 79174 186134 114618
rect 185514 78618 185546 79174
rect 186102 78618 186134 79174
rect 185514 43174 186134 78618
rect 185514 42618 185546 43174
rect 186102 42618 186134 43174
rect 185514 7174 186134 42618
rect 185514 6618 185546 7174
rect 186102 6618 186134 7174
rect 185514 -2266 186134 6618
rect 185514 -2822 185546 -2266
rect 186102 -2822 186134 -2266
rect 185514 -3814 186134 -2822
rect 189234 694894 189854 708122
rect 189234 694338 189266 694894
rect 189822 694338 189854 694894
rect 189234 658894 189854 694338
rect 189234 658338 189266 658894
rect 189822 658338 189854 658894
rect 189234 622894 189854 658338
rect 189234 622338 189266 622894
rect 189822 622338 189854 622894
rect 189234 586894 189854 622338
rect 189234 586338 189266 586894
rect 189822 586338 189854 586894
rect 189234 550894 189854 586338
rect 189234 550338 189266 550894
rect 189822 550338 189854 550894
rect 189234 514894 189854 550338
rect 189234 514338 189266 514894
rect 189822 514338 189854 514894
rect 189234 478894 189854 514338
rect 189234 478338 189266 478894
rect 189822 478338 189854 478894
rect 189234 442894 189854 478338
rect 189234 442338 189266 442894
rect 189822 442338 189854 442894
rect 189234 406894 189854 442338
rect 189234 406338 189266 406894
rect 189822 406338 189854 406894
rect 189234 370894 189854 406338
rect 189234 370338 189266 370894
rect 189822 370338 189854 370894
rect 189234 334894 189854 370338
rect 189234 334338 189266 334894
rect 189822 334338 189854 334894
rect 189234 298894 189854 334338
rect 189234 298338 189266 298894
rect 189822 298338 189854 298894
rect 189234 262894 189854 298338
rect 189234 262338 189266 262894
rect 189822 262338 189854 262894
rect 189234 226894 189854 262338
rect 189234 226338 189266 226894
rect 189822 226338 189854 226894
rect 189234 190894 189854 226338
rect 189234 190338 189266 190894
rect 189822 190338 189854 190894
rect 189234 154894 189854 190338
rect 189234 154338 189266 154894
rect 189822 154338 189854 154894
rect 189234 118894 189854 154338
rect 189234 118338 189266 118894
rect 189822 118338 189854 118894
rect 189234 82894 189854 118338
rect 189234 82338 189266 82894
rect 189822 82338 189854 82894
rect 189234 46894 189854 82338
rect 189234 46338 189266 46894
rect 189822 46338 189854 46894
rect 189234 10894 189854 46338
rect 189234 10338 189266 10894
rect 189822 10338 189854 10894
rect 189234 -4186 189854 10338
rect 189234 -4742 189266 -4186
rect 189822 -4742 189854 -4186
rect 189234 -5734 189854 -4742
rect 192954 698614 193574 710042
rect 210954 711558 211574 711590
rect 210954 711002 210986 711558
rect 211542 711002 211574 711558
rect 207234 709638 207854 709670
rect 207234 709082 207266 709638
rect 207822 709082 207854 709638
rect 203514 707718 204134 707750
rect 203514 707162 203546 707718
rect 204102 707162 204134 707718
rect 192954 698058 192986 698614
rect 193542 698058 193574 698614
rect 192954 662614 193574 698058
rect 192954 662058 192986 662614
rect 193542 662058 193574 662614
rect 192954 626614 193574 662058
rect 192954 626058 192986 626614
rect 193542 626058 193574 626614
rect 192954 590614 193574 626058
rect 192954 590058 192986 590614
rect 193542 590058 193574 590614
rect 192954 554614 193574 590058
rect 192954 554058 192986 554614
rect 193542 554058 193574 554614
rect 192954 518614 193574 554058
rect 192954 518058 192986 518614
rect 193542 518058 193574 518614
rect 192954 482614 193574 518058
rect 192954 482058 192986 482614
rect 193542 482058 193574 482614
rect 192954 446614 193574 482058
rect 192954 446058 192986 446614
rect 193542 446058 193574 446614
rect 192954 410614 193574 446058
rect 192954 410058 192986 410614
rect 193542 410058 193574 410614
rect 192954 374614 193574 410058
rect 192954 374058 192986 374614
rect 193542 374058 193574 374614
rect 192954 338614 193574 374058
rect 192954 338058 192986 338614
rect 193542 338058 193574 338614
rect 192954 302614 193574 338058
rect 192954 302058 192986 302614
rect 193542 302058 193574 302614
rect 192954 266614 193574 302058
rect 192954 266058 192986 266614
rect 193542 266058 193574 266614
rect 192954 230614 193574 266058
rect 192954 230058 192986 230614
rect 193542 230058 193574 230614
rect 192954 194614 193574 230058
rect 192954 194058 192986 194614
rect 193542 194058 193574 194614
rect 192954 158614 193574 194058
rect 192954 158058 192986 158614
rect 193542 158058 193574 158614
rect 192954 122614 193574 158058
rect 192954 122058 192986 122614
rect 193542 122058 193574 122614
rect 192954 86614 193574 122058
rect 192954 86058 192986 86614
rect 193542 86058 193574 86614
rect 192954 50614 193574 86058
rect 192954 50058 192986 50614
rect 193542 50058 193574 50614
rect 192954 14614 193574 50058
rect 192954 14058 192986 14614
rect 193542 14058 193574 14614
rect 174954 -7622 174986 -7066
rect 175542 -7622 175574 -7066
rect 174954 -7654 175574 -7622
rect 192954 -6106 193574 14058
rect 199794 705798 200414 705830
rect 199794 705242 199826 705798
rect 200382 705242 200414 705798
rect 199794 669454 200414 705242
rect 199794 668898 199826 669454
rect 200382 668898 200414 669454
rect 199794 633454 200414 668898
rect 199794 632898 199826 633454
rect 200382 632898 200414 633454
rect 199794 597454 200414 632898
rect 199794 596898 199826 597454
rect 200382 596898 200414 597454
rect 199794 561454 200414 596898
rect 199794 560898 199826 561454
rect 200382 560898 200414 561454
rect 199794 525454 200414 560898
rect 199794 524898 199826 525454
rect 200382 524898 200414 525454
rect 199794 489454 200414 524898
rect 199794 488898 199826 489454
rect 200382 488898 200414 489454
rect 199794 453454 200414 488898
rect 199794 452898 199826 453454
rect 200382 452898 200414 453454
rect 199794 417454 200414 452898
rect 199794 416898 199826 417454
rect 200382 416898 200414 417454
rect 199794 381454 200414 416898
rect 199794 380898 199826 381454
rect 200382 380898 200414 381454
rect 199794 345454 200414 380898
rect 199794 344898 199826 345454
rect 200382 344898 200414 345454
rect 199794 309454 200414 344898
rect 199794 308898 199826 309454
rect 200382 308898 200414 309454
rect 199794 273454 200414 308898
rect 199794 272898 199826 273454
rect 200382 272898 200414 273454
rect 199794 237454 200414 272898
rect 199794 236898 199826 237454
rect 200382 236898 200414 237454
rect 199794 201454 200414 236898
rect 199794 200898 199826 201454
rect 200382 200898 200414 201454
rect 199794 165454 200414 200898
rect 199794 164898 199826 165454
rect 200382 164898 200414 165454
rect 199794 129454 200414 164898
rect 199794 128898 199826 129454
rect 200382 128898 200414 129454
rect 199794 93454 200414 128898
rect 199794 92898 199826 93454
rect 200382 92898 200414 93454
rect 199794 57454 200414 92898
rect 199794 56898 199826 57454
rect 200382 56898 200414 57454
rect 199794 21454 200414 56898
rect 199794 20898 199826 21454
rect 200382 20898 200414 21454
rect 199794 -1306 200414 20898
rect 199794 -1862 199826 -1306
rect 200382 -1862 200414 -1306
rect 199794 -1894 200414 -1862
rect 203514 673174 204134 707162
rect 203514 672618 203546 673174
rect 204102 672618 204134 673174
rect 203514 637174 204134 672618
rect 203514 636618 203546 637174
rect 204102 636618 204134 637174
rect 203514 601174 204134 636618
rect 203514 600618 203546 601174
rect 204102 600618 204134 601174
rect 203514 565174 204134 600618
rect 203514 564618 203546 565174
rect 204102 564618 204134 565174
rect 203514 529174 204134 564618
rect 203514 528618 203546 529174
rect 204102 528618 204134 529174
rect 203514 493174 204134 528618
rect 203514 492618 203546 493174
rect 204102 492618 204134 493174
rect 203514 457174 204134 492618
rect 203514 456618 203546 457174
rect 204102 456618 204134 457174
rect 203514 421174 204134 456618
rect 203514 420618 203546 421174
rect 204102 420618 204134 421174
rect 203514 385174 204134 420618
rect 203514 384618 203546 385174
rect 204102 384618 204134 385174
rect 203514 349174 204134 384618
rect 203514 348618 203546 349174
rect 204102 348618 204134 349174
rect 203514 313174 204134 348618
rect 203514 312618 203546 313174
rect 204102 312618 204134 313174
rect 203514 277174 204134 312618
rect 203514 276618 203546 277174
rect 204102 276618 204134 277174
rect 203514 241174 204134 276618
rect 203514 240618 203546 241174
rect 204102 240618 204134 241174
rect 203514 205174 204134 240618
rect 203514 204618 203546 205174
rect 204102 204618 204134 205174
rect 203514 169174 204134 204618
rect 203514 168618 203546 169174
rect 204102 168618 204134 169174
rect 203514 133174 204134 168618
rect 203514 132618 203546 133174
rect 204102 132618 204134 133174
rect 203514 97174 204134 132618
rect 203514 96618 203546 97174
rect 204102 96618 204134 97174
rect 203514 61174 204134 96618
rect 203514 60618 203546 61174
rect 204102 60618 204134 61174
rect 203514 25174 204134 60618
rect 203514 24618 203546 25174
rect 204102 24618 204134 25174
rect 203514 -3226 204134 24618
rect 203514 -3782 203546 -3226
rect 204102 -3782 204134 -3226
rect 203514 -3814 204134 -3782
rect 207234 676894 207854 709082
rect 207234 676338 207266 676894
rect 207822 676338 207854 676894
rect 207234 640894 207854 676338
rect 207234 640338 207266 640894
rect 207822 640338 207854 640894
rect 207234 604894 207854 640338
rect 207234 604338 207266 604894
rect 207822 604338 207854 604894
rect 207234 568894 207854 604338
rect 207234 568338 207266 568894
rect 207822 568338 207854 568894
rect 207234 532894 207854 568338
rect 207234 532338 207266 532894
rect 207822 532338 207854 532894
rect 207234 496894 207854 532338
rect 207234 496338 207266 496894
rect 207822 496338 207854 496894
rect 207234 460894 207854 496338
rect 207234 460338 207266 460894
rect 207822 460338 207854 460894
rect 207234 424894 207854 460338
rect 207234 424338 207266 424894
rect 207822 424338 207854 424894
rect 207234 388894 207854 424338
rect 207234 388338 207266 388894
rect 207822 388338 207854 388894
rect 207234 352894 207854 388338
rect 207234 352338 207266 352894
rect 207822 352338 207854 352894
rect 207234 316894 207854 352338
rect 207234 316338 207266 316894
rect 207822 316338 207854 316894
rect 207234 280894 207854 316338
rect 207234 280338 207266 280894
rect 207822 280338 207854 280894
rect 207234 244894 207854 280338
rect 207234 244338 207266 244894
rect 207822 244338 207854 244894
rect 207234 208894 207854 244338
rect 207234 208338 207266 208894
rect 207822 208338 207854 208894
rect 207234 172894 207854 208338
rect 207234 172338 207266 172894
rect 207822 172338 207854 172894
rect 207234 136894 207854 172338
rect 207234 136338 207266 136894
rect 207822 136338 207854 136894
rect 207234 100894 207854 136338
rect 207234 100338 207266 100894
rect 207822 100338 207854 100894
rect 207234 64894 207854 100338
rect 207234 64338 207266 64894
rect 207822 64338 207854 64894
rect 207234 28894 207854 64338
rect 207234 28338 207266 28894
rect 207822 28338 207854 28894
rect 207234 -5146 207854 28338
rect 207234 -5702 207266 -5146
rect 207822 -5702 207854 -5146
rect 207234 -5734 207854 -5702
rect 210954 680614 211574 711002
rect 228954 710598 229574 711590
rect 228954 710042 228986 710598
rect 229542 710042 229574 710598
rect 225234 708678 225854 709670
rect 225234 708122 225266 708678
rect 225822 708122 225854 708678
rect 221514 706758 222134 707750
rect 221514 706202 221546 706758
rect 222102 706202 222134 706758
rect 210954 680058 210986 680614
rect 211542 680058 211574 680614
rect 210954 644614 211574 680058
rect 210954 644058 210986 644614
rect 211542 644058 211574 644614
rect 210954 608614 211574 644058
rect 210954 608058 210986 608614
rect 211542 608058 211574 608614
rect 210954 572614 211574 608058
rect 210954 572058 210986 572614
rect 211542 572058 211574 572614
rect 210954 536614 211574 572058
rect 210954 536058 210986 536614
rect 211542 536058 211574 536614
rect 210954 500614 211574 536058
rect 210954 500058 210986 500614
rect 211542 500058 211574 500614
rect 210954 464614 211574 500058
rect 210954 464058 210986 464614
rect 211542 464058 211574 464614
rect 210954 428614 211574 464058
rect 210954 428058 210986 428614
rect 211542 428058 211574 428614
rect 210954 392614 211574 428058
rect 210954 392058 210986 392614
rect 211542 392058 211574 392614
rect 210954 356614 211574 392058
rect 210954 356058 210986 356614
rect 211542 356058 211574 356614
rect 210954 320614 211574 356058
rect 210954 320058 210986 320614
rect 211542 320058 211574 320614
rect 210954 284614 211574 320058
rect 210954 284058 210986 284614
rect 211542 284058 211574 284614
rect 210954 248614 211574 284058
rect 210954 248058 210986 248614
rect 211542 248058 211574 248614
rect 210954 212614 211574 248058
rect 210954 212058 210986 212614
rect 211542 212058 211574 212614
rect 210954 176614 211574 212058
rect 210954 176058 210986 176614
rect 211542 176058 211574 176614
rect 210954 140614 211574 176058
rect 210954 140058 210986 140614
rect 211542 140058 211574 140614
rect 210954 104614 211574 140058
rect 210954 104058 210986 104614
rect 211542 104058 211574 104614
rect 210954 68614 211574 104058
rect 210954 68058 210986 68614
rect 211542 68058 211574 68614
rect 210954 32614 211574 68058
rect 210954 32058 210986 32614
rect 211542 32058 211574 32614
rect 192954 -6662 192986 -6106
rect 193542 -6662 193574 -6106
rect 192954 -7654 193574 -6662
rect 210954 -7066 211574 32058
rect 217794 704838 218414 705830
rect 217794 704282 217826 704838
rect 218382 704282 218414 704838
rect 217794 687454 218414 704282
rect 217794 686898 217826 687454
rect 218382 686898 218414 687454
rect 217794 651454 218414 686898
rect 217794 650898 217826 651454
rect 218382 650898 218414 651454
rect 217794 615454 218414 650898
rect 217794 614898 217826 615454
rect 218382 614898 218414 615454
rect 217794 579454 218414 614898
rect 217794 578898 217826 579454
rect 218382 578898 218414 579454
rect 217794 543454 218414 578898
rect 217794 542898 217826 543454
rect 218382 542898 218414 543454
rect 217794 507454 218414 542898
rect 217794 506898 217826 507454
rect 218382 506898 218414 507454
rect 217794 471454 218414 506898
rect 217794 470898 217826 471454
rect 218382 470898 218414 471454
rect 217794 435454 218414 470898
rect 217794 434898 217826 435454
rect 218382 434898 218414 435454
rect 217794 399454 218414 434898
rect 217794 398898 217826 399454
rect 218382 398898 218414 399454
rect 217794 363454 218414 398898
rect 217794 362898 217826 363454
rect 218382 362898 218414 363454
rect 217794 327454 218414 362898
rect 217794 326898 217826 327454
rect 218382 326898 218414 327454
rect 217794 291454 218414 326898
rect 217794 290898 217826 291454
rect 218382 290898 218414 291454
rect 217794 255454 218414 290898
rect 217794 254898 217826 255454
rect 218382 254898 218414 255454
rect 217794 219454 218414 254898
rect 217794 218898 217826 219454
rect 218382 218898 218414 219454
rect 217794 183454 218414 218898
rect 217794 182898 217826 183454
rect 218382 182898 218414 183454
rect 217794 147454 218414 182898
rect 217794 146898 217826 147454
rect 218382 146898 218414 147454
rect 217794 111454 218414 146898
rect 217794 110898 217826 111454
rect 218382 110898 218414 111454
rect 217794 75454 218414 110898
rect 217794 74898 217826 75454
rect 218382 74898 218414 75454
rect 217794 39454 218414 74898
rect 217794 38898 217826 39454
rect 218382 38898 218414 39454
rect 217794 3454 218414 38898
rect 217794 2898 217826 3454
rect 218382 2898 218414 3454
rect 217794 -346 218414 2898
rect 217794 -902 217826 -346
rect 218382 -902 218414 -346
rect 217794 -1894 218414 -902
rect 221514 691174 222134 706202
rect 221514 690618 221546 691174
rect 222102 690618 222134 691174
rect 221514 655174 222134 690618
rect 221514 654618 221546 655174
rect 222102 654618 222134 655174
rect 221514 619174 222134 654618
rect 221514 618618 221546 619174
rect 222102 618618 222134 619174
rect 221514 583174 222134 618618
rect 221514 582618 221546 583174
rect 222102 582618 222134 583174
rect 221514 547174 222134 582618
rect 221514 546618 221546 547174
rect 222102 546618 222134 547174
rect 221514 511174 222134 546618
rect 221514 510618 221546 511174
rect 222102 510618 222134 511174
rect 221514 475174 222134 510618
rect 221514 474618 221546 475174
rect 222102 474618 222134 475174
rect 221514 439174 222134 474618
rect 221514 438618 221546 439174
rect 222102 438618 222134 439174
rect 221514 403174 222134 438618
rect 221514 402618 221546 403174
rect 222102 402618 222134 403174
rect 221514 367174 222134 402618
rect 221514 366618 221546 367174
rect 222102 366618 222134 367174
rect 221514 331174 222134 366618
rect 221514 330618 221546 331174
rect 222102 330618 222134 331174
rect 221514 295174 222134 330618
rect 221514 294618 221546 295174
rect 222102 294618 222134 295174
rect 221514 259174 222134 294618
rect 221514 258618 221546 259174
rect 222102 258618 222134 259174
rect 221514 223174 222134 258618
rect 221514 222618 221546 223174
rect 222102 222618 222134 223174
rect 221514 187174 222134 222618
rect 221514 186618 221546 187174
rect 222102 186618 222134 187174
rect 221514 151174 222134 186618
rect 221514 150618 221546 151174
rect 222102 150618 222134 151174
rect 221514 115174 222134 150618
rect 221514 114618 221546 115174
rect 222102 114618 222134 115174
rect 221514 79174 222134 114618
rect 221514 78618 221546 79174
rect 222102 78618 222134 79174
rect 221514 43174 222134 78618
rect 221514 42618 221546 43174
rect 222102 42618 222134 43174
rect 221514 7174 222134 42618
rect 221514 6618 221546 7174
rect 222102 6618 222134 7174
rect 221514 -2266 222134 6618
rect 221514 -2822 221546 -2266
rect 222102 -2822 222134 -2266
rect 221514 -3814 222134 -2822
rect 225234 694894 225854 708122
rect 225234 694338 225266 694894
rect 225822 694338 225854 694894
rect 225234 658894 225854 694338
rect 225234 658338 225266 658894
rect 225822 658338 225854 658894
rect 225234 622894 225854 658338
rect 225234 622338 225266 622894
rect 225822 622338 225854 622894
rect 225234 586894 225854 622338
rect 225234 586338 225266 586894
rect 225822 586338 225854 586894
rect 225234 550894 225854 586338
rect 225234 550338 225266 550894
rect 225822 550338 225854 550894
rect 225234 514894 225854 550338
rect 225234 514338 225266 514894
rect 225822 514338 225854 514894
rect 225234 478894 225854 514338
rect 225234 478338 225266 478894
rect 225822 478338 225854 478894
rect 225234 442894 225854 478338
rect 225234 442338 225266 442894
rect 225822 442338 225854 442894
rect 225234 406894 225854 442338
rect 225234 406338 225266 406894
rect 225822 406338 225854 406894
rect 225234 370894 225854 406338
rect 225234 370338 225266 370894
rect 225822 370338 225854 370894
rect 225234 334894 225854 370338
rect 225234 334338 225266 334894
rect 225822 334338 225854 334894
rect 225234 298894 225854 334338
rect 225234 298338 225266 298894
rect 225822 298338 225854 298894
rect 225234 262894 225854 298338
rect 225234 262338 225266 262894
rect 225822 262338 225854 262894
rect 225234 226894 225854 262338
rect 225234 226338 225266 226894
rect 225822 226338 225854 226894
rect 225234 190894 225854 226338
rect 225234 190338 225266 190894
rect 225822 190338 225854 190894
rect 225234 154894 225854 190338
rect 225234 154338 225266 154894
rect 225822 154338 225854 154894
rect 225234 118894 225854 154338
rect 225234 118338 225266 118894
rect 225822 118338 225854 118894
rect 225234 82894 225854 118338
rect 225234 82338 225266 82894
rect 225822 82338 225854 82894
rect 225234 46894 225854 82338
rect 225234 46338 225266 46894
rect 225822 46338 225854 46894
rect 225234 10894 225854 46338
rect 225234 10338 225266 10894
rect 225822 10338 225854 10894
rect 225234 -4186 225854 10338
rect 225234 -4742 225266 -4186
rect 225822 -4742 225854 -4186
rect 225234 -5734 225854 -4742
rect 228954 698614 229574 710042
rect 246954 711558 247574 711590
rect 246954 711002 246986 711558
rect 247542 711002 247574 711558
rect 243234 709638 243854 709670
rect 243234 709082 243266 709638
rect 243822 709082 243854 709638
rect 239514 707718 240134 707750
rect 239514 707162 239546 707718
rect 240102 707162 240134 707718
rect 228954 698058 228986 698614
rect 229542 698058 229574 698614
rect 228954 662614 229574 698058
rect 228954 662058 228986 662614
rect 229542 662058 229574 662614
rect 228954 626614 229574 662058
rect 228954 626058 228986 626614
rect 229542 626058 229574 626614
rect 228954 590614 229574 626058
rect 228954 590058 228986 590614
rect 229542 590058 229574 590614
rect 228954 554614 229574 590058
rect 228954 554058 228986 554614
rect 229542 554058 229574 554614
rect 228954 518614 229574 554058
rect 228954 518058 228986 518614
rect 229542 518058 229574 518614
rect 228954 482614 229574 518058
rect 235794 705798 236414 705830
rect 235794 705242 235826 705798
rect 236382 705242 236414 705798
rect 235794 669454 236414 705242
rect 235794 668898 235826 669454
rect 236382 668898 236414 669454
rect 235794 633454 236414 668898
rect 235794 632898 235826 633454
rect 236382 632898 236414 633454
rect 235794 597454 236414 632898
rect 235794 596898 235826 597454
rect 236382 596898 236414 597454
rect 235794 561454 236414 596898
rect 235794 560898 235826 561454
rect 236382 560898 236414 561454
rect 235794 525454 236414 560898
rect 235794 524898 235826 525454
rect 236382 524898 236414 525454
rect 235794 489603 236414 524898
rect 239514 673174 240134 707162
rect 239514 672618 239546 673174
rect 240102 672618 240134 673174
rect 239514 637174 240134 672618
rect 239514 636618 239546 637174
rect 240102 636618 240134 637174
rect 239514 601174 240134 636618
rect 239514 600618 239546 601174
rect 240102 600618 240134 601174
rect 239514 565174 240134 600618
rect 239514 564618 239546 565174
rect 240102 564618 240134 565174
rect 239514 529174 240134 564618
rect 239514 528618 239546 529174
rect 240102 528618 240134 529174
rect 239514 493174 240134 528618
rect 239514 492618 239546 493174
rect 240102 492618 240134 493174
rect 239514 489603 240134 492618
rect 243234 676894 243854 709082
rect 243234 676338 243266 676894
rect 243822 676338 243854 676894
rect 243234 640894 243854 676338
rect 243234 640338 243266 640894
rect 243822 640338 243854 640894
rect 243234 604894 243854 640338
rect 243234 604338 243266 604894
rect 243822 604338 243854 604894
rect 243234 568894 243854 604338
rect 243234 568338 243266 568894
rect 243822 568338 243854 568894
rect 243234 532894 243854 568338
rect 243234 532338 243266 532894
rect 243822 532338 243854 532894
rect 243234 496894 243854 532338
rect 243234 496338 243266 496894
rect 243822 496338 243854 496894
rect 243234 489603 243854 496338
rect 246954 680614 247574 711002
rect 264954 710598 265574 711590
rect 264954 710042 264986 710598
rect 265542 710042 265574 710598
rect 261234 708678 261854 709670
rect 261234 708122 261266 708678
rect 261822 708122 261854 708678
rect 257514 706758 258134 707750
rect 257514 706202 257546 706758
rect 258102 706202 258134 706758
rect 246954 680058 246986 680614
rect 247542 680058 247574 680614
rect 246954 644614 247574 680058
rect 246954 644058 246986 644614
rect 247542 644058 247574 644614
rect 246954 608614 247574 644058
rect 246954 608058 246986 608614
rect 247542 608058 247574 608614
rect 246954 572614 247574 608058
rect 246954 572058 246986 572614
rect 247542 572058 247574 572614
rect 246954 536614 247574 572058
rect 246954 536058 246986 536614
rect 247542 536058 247574 536614
rect 246954 500614 247574 536058
rect 246954 500058 246986 500614
rect 247542 500058 247574 500614
rect 246954 489603 247574 500058
rect 253794 704838 254414 705830
rect 253794 704282 253826 704838
rect 254382 704282 254414 704838
rect 253794 687454 254414 704282
rect 253794 686898 253826 687454
rect 254382 686898 254414 687454
rect 253794 651454 254414 686898
rect 253794 650898 253826 651454
rect 254382 650898 254414 651454
rect 253794 615454 254414 650898
rect 253794 614898 253826 615454
rect 254382 614898 254414 615454
rect 253794 579454 254414 614898
rect 253794 578898 253826 579454
rect 254382 578898 254414 579454
rect 253794 543454 254414 578898
rect 253794 542898 253826 543454
rect 254382 542898 254414 543454
rect 253794 507454 254414 542898
rect 253794 506898 253826 507454
rect 254382 506898 254414 507454
rect 253794 489603 254414 506898
rect 257514 691174 258134 706202
rect 257514 690618 257546 691174
rect 258102 690618 258134 691174
rect 257514 655174 258134 690618
rect 257514 654618 257546 655174
rect 258102 654618 258134 655174
rect 257514 619174 258134 654618
rect 257514 618618 257546 619174
rect 258102 618618 258134 619174
rect 257514 583174 258134 618618
rect 257514 582618 257546 583174
rect 258102 582618 258134 583174
rect 257514 547174 258134 582618
rect 257514 546618 257546 547174
rect 258102 546618 258134 547174
rect 257514 511174 258134 546618
rect 257514 510618 257546 511174
rect 258102 510618 258134 511174
rect 257514 489603 258134 510618
rect 261234 694894 261854 708122
rect 261234 694338 261266 694894
rect 261822 694338 261854 694894
rect 261234 658894 261854 694338
rect 261234 658338 261266 658894
rect 261822 658338 261854 658894
rect 261234 622894 261854 658338
rect 261234 622338 261266 622894
rect 261822 622338 261854 622894
rect 261234 586894 261854 622338
rect 261234 586338 261266 586894
rect 261822 586338 261854 586894
rect 261234 550894 261854 586338
rect 261234 550338 261266 550894
rect 261822 550338 261854 550894
rect 261234 514894 261854 550338
rect 261234 514338 261266 514894
rect 261822 514338 261854 514894
rect 261234 489603 261854 514338
rect 264954 698614 265574 710042
rect 282954 711558 283574 711590
rect 282954 711002 282986 711558
rect 283542 711002 283574 711558
rect 279234 709638 279854 709670
rect 279234 709082 279266 709638
rect 279822 709082 279854 709638
rect 275514 707718 276134 707750
rect 275514 707162 275546 707718
rect 276102 707162 276134 707718
rect 264954 698058 264986 698614
rect 265542 698058 265574 698614
rect 264954 662614 265574 698058
rect 264954 662058 264986 662614
rect 265542 662058 265574 662614
rect 264954 626614 265574 662058
rect 264954 626058 264986 626614
rect 265542 626058 265574 626614
rect 264954 590614 265574 626058
rect 264954 590058 264986 590614
rect 265542 590058 265574 590614
rect 264954 554614 265574 590058
rect 264954 554058 264986 554614
rect 265542 554058 265574 554614
rect 264954 518614 265574 554058
rect 264954 518058 264986 518614
rect 265542 518058 265574 518614
rect 264954 489603 265574 518058
rect 271794 705798 272414 705830
rect 271794 705242 271826 705798
rect 272382 705242 272414 705798
rect 271794 669454 272414 705242
rect 271794 668898 271826 669454
rect 272382 668898 272414 669454
rect 271794 633454 272414 668898
rect 271794 632898 271826 633454
rect 272382 632898 272414 633454
rect 271794 597454 272414 632898
rect 271794 596898 271826 597454
rect 272382 596898 272414 597454
rect 271794 561454 272414 596898
rect 271794 560898 271826 561454
rect 272382 560898 272414 561454
rect 271794 525454 272414 560898
rect 271794 524898 271826 525454
rect 272382 524898 272414 525454
rect 271794 489603 272414 524898
rect 275514 673174 276134 707162
rect 275514 672618 275546 673174
rect 276102 672618 276134 673174
rect 275514 637174 276134 672618
rect 275514 636618 275546 637174
rect 276102 636618 276134 637174
rect 275514 601174 276134 636618
rect 275514 600618 275546 601174
rect 276102 600618 276134 601174
rect 275514 565174 276134 600618
rect 275514 564618 275546 565174
rect 276102 564618 276134 565174
rect 275514 529174 276134 564618
rect 275514 528618 275546 529174
rect 276102 528618 276134 529174
rect 275514 493174 276134 528618
rect 275514 492618 275546 493174
rect 276102 492618 276134 493174
rect 275514 489603 276134 492618
rect 279234 676894 279854 709082
rect 279234 676338 279266 676894
rect 279822 676338 279854 676894
rect 279234 640894 279854 676338
rect 279234 640338 279266 640894
rect 279822 640338 279854 640894
rect 279234 604894 279854 640338
rect 279234 604338 279266 604894
rect 279822 604338 279854 604894
rect 279234 568894 279854 604338
rect 279234 568338 279266 568894
rect 279822 568338 279854 568894
rect 279234 532894 279854 568338
rect 279234 532338 279266 532894
rect 279822 532338 279854 532894
rect 279234 496894 279854 532338
rect 279234 496338 279266 496894
rect 279822 496338 279854 496894
rect 279234 489603 279854 496338
rect 282954 680614 283574 711002
rect 300954 710598 301574 711590
rect 300954 710042 300986 710598
rect 301542 710042 301574 710598
rect 297234 708678 297854 709670
rect 297234 708122 297266 708678
rect 297822 708122 297854 708678
rect 293514 706758 294134 707750
rect 293514 706202 293546 706758
rect 294102 706202 294134 706758
rect 282954 680058 282986 680614
rect 283542 680058 283574 680614
rect 282954 644614 283574 680058
rect 282954 644058 282986 644614
rect 283542 644058 283574 644614
rect 282954 608614 283574 644058
rect 282954 608058 282986 608614
rect 283542 608058 283574 608614
rect 282954 572614 283574 608058
rect 282954 572058 282986 572614
rect 283542 572058 283574 572614
rect 282954 536614 283574 572058
rect 282954 536058 282986 536614
rect 283542 536058 283574 536614
rect 282954 500614 283574 536058
rect 282954 500058 282986 500614
rect 283542 500058 283574 500614
rect 282954 489603 283574 500058
rect 289794 704838 290414 705830
rect 289794 704282 289826 704838
rect 290382 704282 290414 704838
rect 289794 687454 290414 704282
rect 289794 686898 289826 687454
rect 290382 686898 290414 687454
rect 289794 651454 290414 686898
rect 289794 650898 289826 651454
rect 290382 650898 290414 651454
rect 289794 615454 290414 650898
rect 289794 614898 289826 615454
rect 290382 614898 290414 615454
rect 289794 579454 290414 614898
rect 289794 578898 289826 579454
rect 290382 578898 290414 579454
rect 289794 543454 290414 578898
rect 289794 542898 289826 543454
rect 290382 542898 290414 543454
rect 289794 507454 290414 542898
rect 289794 506898 289826 507454
rect 290382 506898 290414 507454
rect 289794 489603 290414 506898
rect 293514 691174 294134 706202
rect 293514 690618 293546 691174
rect 294102 690618 294134 691174
rect 293514 655174 294134 690618
rect 293514 654618 293546 655174
rect 294102 654618 294134 655174
rect 293514 619174 294134 654618
rect 293514 618618 293546 619174
rect 294102 618618 294134 619174
rect 293514 583174 294134 618618
rect 293514 582618 293546 583174
rect 294102 582618 294134 583174
rect 293514 547174 294134 582618
rect 293514 546618 293546 547174
rect 294102 546618 294134 547174
rect 293514 511174 294134 546618
rect 293514 510618 293546 511174
rect 294102 510618 294134 511174
rect 293514 489603 294134 510618
rect 297234 694894 297854 708122
rect 297234 694338 297266 694894
rect 297822 694338 297854 694894
rect 297234 658894 297854 694338
rect 297234 658338 297266 658894
rect 297822 658338 297854 658894
rect 297234 622894 297854 658338
rect 297234 622338 297266 622894
rect 297822 622338 297854 622894
rect 297234 586894 297854 622338
rect 297234 586338 297266 586894
rect 297822 586338 297854 586894
rect 297234 550894 297854 586338
rect 297234 550338 297266 550894
rect 297822 550338 297854 550894
rect 297234 514894 297854 550338
rect 297234 514338 297266 514894
rect 297822 514338 297854 514894
rect 297234 489603 297854 514338
rect 300954 698614 301574 710042
rect 318954 711558 319574 711590
rect 318954 711002 318986 711558
rect 319542 711002 319574 711558
rect 315234 709638 315854 709670
rect 315234 709082 315266 709638
rect 315822 709082 315854 709638
rect 311514 707718 312134 707750
rect 311514 707162 311546 707718
rect 312102 707162 312134 707718
rect 300954 698058 300986 698614
rect 301542 698058 301574 698614
rect 300954 662614 301574 698058
rect 300954 662058 300986 662614
rect 301542 662058 301574 662614
rect 300954 626614 301574 662058
rect 300954 626058 300986 626614
rect 301542 626058 301574 626614
rect 300954 590614 301574 626058
rect 300954 590058 300986 590614
rect 301542 590058 301574 590614
rect 300954 554614 301574 590058
rect 300954 554058 300986 554614
rect 301542 554058 301574 554614
rect 300954 518614 301574 554058
rect 300954 518058 300986 518614
rect 301542 518058 301574 518614
rect 300954 489603 301574 518058
rect 307794 705798 308414 705830
rect 307794 705242 307826 705798
rect 308382 705242 308414 705798
rect 307794 669454 308414 705242
rect 307794 668898 307826 669454
rect 308382 668898 308414 669454
rect 307794 633454 308414 668898
rect 307794 632898 307826 633454
rect 308382 632898 308414 633454
rect 307794 597454 308414 632898
rect 307794 596898 307826 597454
rect 308382 596898 308414 597454
rect 307794 561454 308414 596898
rect 307794 560898 307826 561454
rect 308382 560898 308414 561454
rect 307794 525454 308414 560898
rect 307794 524898 307826 525454
rect 308382 524898 308414 525454
rect 307794 489603 308414 524898
rect 311514 673174 312134 707162
rect 311514 672618 311546 673174
rect 312102 672618 312134 673174
rect 311514 637174 312134 672618
rect 311514 636618 311546 637174
rect 312102 636618 312134 637174
rect 311514 601174 312134 636618
rect 311514 600618 311546 601174
rect 312102 600618 312134 601174
rect 311514 565174 312134 600618
rect 311514 564618 311546 565174
rect 312102 564618 312134 565174
rect 311514 529174 312134 564618
rect 311514 528618 311546 529174
rect 312102 528618 312134 529174
rect 311514 493174 312134 528618
rect 311514 492618 311546 493174
rect 312102 492618 312134 493174
rect 311514 489603 312134 492618
rect 315234 676894 315854 709082
rect 315234 676338 315266 676894
rect 315822 676338 315854 676894
rect 315234 640894 315854 676338
rect 315234 640338 315266 640894
rect 315822 640338 315854 640894
rect 315234 604894 315854 640338
rect 315234 604338 315266 604894
rect 315822 604338 315854 604894
rect 315234 568894 315854 604338
rect 315234 568338 315266 568894
rect 315822 568338 315854 568894
rect 315234 532894 315854 568338
rect 315234 532338 315266 532894
rect 315822 532338 315854 532894
rect 315234 496894 315854 532338
rect 315234 496338 315266 496894
rect 315822 496338 315854 496894
rect 315234 489603 315854 496338
rect 318954 680614 319574 711002
rect 336954 710598 337574 711590
rect 336954 710042 336986 710598
rect 337542 710042 337574 710598
rect 333234 708678 333854 709670
rect 333234 708122 333266 708678
rect 333822 708122 333854 708678
rect 329514 706758 330134 707750
rect 329514 706202 329546 706758
rect 330102 706202 330134 706758
rect 318954 680058 318986 680614
rect 319542 680058 319574 680614
rect 318954 644614 319574 680058
rect 318954 644058 318986 644614
rect 319542 644058 319574 644614
rect 318954 608614 319574 644058
rect 318954 608058 318986 608614
rect 319542 608058 319574 608614
rect 318954 572614 319574 608058
rect 318954 572058 318986 572614
rect 319542 572058 319574 572614
rect 318954 536614 319574 572058
rect 318954 536058 318986 536614
rect 319542 536058 319574 536614
rect 318954 500614 319574 536058
rect 318954 500058 318986 500614
rect 319542 500058 319574 500614
rect 318954 489603 319574 500058
rect 325794 704838 326414 705830
rect 325794 704282 325826 704838
rect 326382 704282 326414 704838
rect 325794 687454 326414 704282
rect 325794 686898 325826 687454
rect 326382 686898 326414 687454
rect 325794 651454 326414 686898
rect 325794 650898 325826 651454
rect 326382 650898 326414 651454
rect 325794 615454 326414 650898
rect 325794 614898 325826 615454
rect 326382 614898 326414 615454
rect 325794 579454 326414 614898
rect 325794 578898 325826 579454
rect 326382 578898 326414 579454
rect 325794 543454 326414 578898
rect 325794 542898 325826 543454
rect 326382 542898 326414 543454
rect 325794 507454 326414 542898
rect 325794 506898 325826 507454
rect 326382 506898 326414 507454
rect 325794 489603 326414 506898
rect 329514 691174 330134 706202
rect 329514 690618 329546 691174
rect 330102 690618 330134 691174
rect 329514 655174 330134 690618
rect 329514 654618 329546 655174
rect 330102 654618 330134 655174
rect 329514 619174 330134 654618
rect 329514 618618 329546 619174
rect 330102 618618 330134 619174
rect 329514 583174 330134 618618
rect 329514 582618 329546 583174
rect 330102 582618 330134 583174
rect 329514 547174 330134 582618
rect 329514 546618 329546 547174
rect 330102 546618 330134 547174
rect 329514 511174 330134 546618
rect 329514 510618 329546 511174
rect 330102 510618 330134 511174
rect 329514 489603 330134 510618
rect 333234 694894 333854 708122
rect 333234 694338 333266 694894
rect 333822 694338 333854 694894
rect 333234 658894 333854 694338
rect 333234 658338 333266 658894
rect 333822 658338 333854 658894
rect 333234 622894 333854 658338
rect 333234 622338 333266 622894
rect 333822 622338 333854 622894
rect 333234 586894 333854 622338
rect 333234 586338 333266 586894
rect 333822 586338 333854 586894
rect 333234 550894 333854 586338
rect 333234 550338 333266 550894
rect 333822 550338 333854 550894
rect 333234 514894 333854 550338
rect 333234 514338 333266 514894
rect 333822 514338 333854 514894
rect 333234 489603 333854 514338
rect 336954 698614 337574 710042
rect 354954 711558 355574 711590
rect 354954 711002 354986 711558
rect 355542 711002 355574 711558
rect 351234 709638 351854 709670
rect 351234 709082 351266 709638
rect 351822 709082 351854 709638
rect 347514 707718 348134 707750
rect 347514 707162 347546 707718
rect 348102 707162 348134 707718
rect 336954 698058 336986 698614
rect 337542 698058 337574 698614
rect 336954 662614 337574 698058
rect 336954 662058 336986 662614
rect 337542 662058 337574 662614
rect 336954 626614 337574 662058
rect 336954 626058 336986 626614
rect 337542 626058 337574 626614
rect 336954 590614 337574 626058
rect 336954 590058 336986 590614
rect 337542 590058 337574 590614
rect 336954 554614 337574 590058
rect 336954 554058 336986 554614
rect 337542 554058 337574 554614
rect 336954 518614 337574 554058
rect 336954 518058 336986 518614
rect 337542 518058 337574 518614
rect 336954 489603 337574 518058
rect 343794 705798 344414 705830
rect 343794 705242 343826 705798
rect 344382 705242 344414 705798
rect 343794 669454 344414 705242
rect 343794 668898 343826 669454
rect 344382 668898 344414 669454
rect 343794 633454 344414 668898
rect 343794 632898 343826 633454
rect 344382 632898 344414 633454
rect 343794 597454 344414 632898
rect 343794 596898 343826 597454
rect 344382 596898 344414 597454
rect 343794 561454 344414 596898
rect 343794 560898 343826 561454
rect 344382 560898 344414 561454
rect 343794 525454 344414 560898
rect 343794 524898 343826 525454
rect 344382 524898 344414 525454
rect 343794 489603 344414 524898
rect 347514 673174 348134 707162
rect 347514 672618 347546 673174
rect 348102 672618 348134 673174
rect 347514 637174 348134 672618
rect 347514 636618 347546 637174
rect 348102 636618 348134 637174
rect 347514 601174 348134 636618
rect 347514 600618 347546 601174
rect 348102 600618 348134 601174
rect 347514 565174 348134 600618
rect 347514 564618 347546 565174
rect 348102 564618 348134 565174
rect 347514 529174 348134 564618
rect 347514 528618 347546 529174
rect 348102 528618 348134 529174
rect 347514 493174 348134 528618
rect 347514 492618 347546 493174
rect 348102 492618 348134 493174
rect 347514 489603 348134 492618
rect 351234 676894 351854 709082
rect 351234 676338 351266 676894
rect 351822 676338 351854 676894
rect 351234 640894 351854 676338
rect 351234 640338 351266 640894
rect 351822 640338 351854 640894
rect 351234 604894 351854 640338
rect 351234 604338 351266 604894
rect 351822 604338 351854 604894
rect 351234 568894 351854 604338
rect 351234 568338 351266 568894
rect 351822 568338 351854 568894
rect 351234 532894 351854 568338
rect 351234 532338 351266 532894
rect 351822 532338 351854 532894
rect 351234 496894 351854 532338
rect 351234 496338 351266 496894
rect 351822 496338 351854 496894
rect 351234 489603 351854 496338
rect 354954 680614 355574 711002
rect 372954 710598 373574 711590
rect 372954 710042 372986 710598
rect 373542 710042 373574 710598
rect 369234 708678 369854 709670
rect 369234 708122 369266 708678
rect 369822 708122 369854 708678
rect 365514 706758 366134 707750
rect 365514 706202 365546 706758
rect 366102 706202 366134 706758
rect 354954 680058 354986 680614
rect 355542 680058 355574 680614
rect 354954 644614 355574 680058
rect 354954 644058 354986 644614
rect 355542 644058 355574 644614
rect 354954 608614 355574 644058
rect 354954 608058 354986 608614
rect 355542 608058 355574 608614
rect 354954 572614 355574 608058
rect 354954 572058 354986 572614
rect 355542 572058 355574 572614
rect 354954 536614 355574 572058
rect 354954 536058 354986 536614
rect 355542 536058 355574 536614
rect 354954 500614 355574 536058
rect 354954 500058 354986 500614
rect 355542 500058 355574 500614
rect 354954 489603 355574 500058
rect 361794 704838 362414 705830
rect 361794 704282 361826 704838
rect 362382 704282 362414 704838
rect 361794 687454 362414 704282
rect 361794 686898 361826 687454
rect 362382 686898 362414 687454
rect 361794 651454 362414 686898
rect 361794 650898 361826 651454
rect 362382 650898 362414 651454
rect 361794 615454 362414 650898
rect 361794 614898 361826 615454
rect 362382 614898 362414 615454
rect 361794 579454 362414 614898
rect 361794 578898 361826 579454
rect 362382 578898 362414 579454
rect 361794 543454 362414 578898
rect 361794 542898 361826 543454
rect 362382 542898 362414 543454
rect 361794 507454 362414 542898
rect 361794 506898 361826 507454
rect 362382 506898 362414 507454
rect 361794 489603 362414 506898
rect 365514 691174 366134 706202
rect 365514 690618 365546 691174
rect 366102 690618 366134 691174
rect 365514 655174 366134 690618
rect 365514 654618 365546 655174
rect 366102 654618 366134 655174
rect 365514 619174 366134 654618
rect 365514 618618 365546 619174
rect 366102 618618 366134 619174
rect 365514 583174 366134 618618
rect 365514 582618 365546 583174
rect 366102 582618 366134 583174
rect 365514 547174 366134 582618
rect 365514 546618 365546 547174
rect 366102 546618 366134 547174
rect 365514 511174 366134 546618
rect 365514 510618 365546 511174
rect 366102 510618 366134 511174
rect 365514 489603 366134 510618
rect 369234 694894 369854 708122
rect 369234 694338 369266 694894
rect 369822 694338 369854 694894
rect 369234 658894 369854 694338
rect 369234 658338 369266 658894
rect 369822 658338 369854 658894
rect 369234 622894 369854 658338
rect 369234 622338 369266 622894
rect 369822 622338 369854 622894
rect 369234 586894 369854 622338
rect 369234 586338 369266 586894
rect 369822 586338 369854 586894
rect 369234 550894 369854 586338
rect 369234 550338 369266 550894
rect 369822 550338 369854 550894
rect 369234 514894 369854 550338
rect 369234 514338 369266 514894
rect 369822 514338 369854 514894
rect 369234 489603 369854 514338
rect 372954 698614 373574 710042
rect 390954 711558 391574 711590
rect 390954 711002 390986 711558
rect 391542 711002 391574 711558
rect 387234 709638 387854 709670
rect 387234 709082 387266 709638
rect 387822 709082 387854 709638
rect 383514 707718 384134 707750
rect 383514 707162 383546 707718
rect 384102 707162 384134 707718
rect 372954 698058 372986 698614
rect 373542 698058 373574 698614
rect 372954 662614 373574 698058
rect 372954 662058 372986 662614
rect 373542 662058 373574 662614
rect 372954 626614 373574 662058
rect 372954 626058 372986 626614
rect 373542 626058 373574 626614
rect 372954 590614 373574 626058
rect 372954 590058 372986 590614
rect 373542 590058 373574 590614
rect 372954 554614 373574 590058
rect 372954 554058 372986 554614
rect 373542 554058 373574 554614
rect 372954 518614 373574 554058
rect 372954 518058 372986 518614
rect 373542 518058 373574 518614
rect 372954 489603 373574 518058
rect 379794 705798 380414 705830
rect 379794 705242 379826 705798
rect 380382 705242 380414 705798
rect 379794 669454 380414 705242
rect 379794 668898 379826 669454
rect 380382 668898 380414 669454
rect 379794 633454 380414 668898
rect 379794 632898 379826 633454
rect 380382 632898 380414 633454
rect 379794 597454 380414 632898
rect 379794 596898 379826 597454
rect 380382 596898 380414 597454
rect 379794 561454 380414 596898
rect 379794 560898 379826 561454
rect 380382 560898 380414 561454
rect 379794 525454 380414 560898
rect 379794 524898 379826 525454
rect 380382 524898 380414 525454
rect 379794 489603 380414 524898
rect 383514 673174 384134 707162
rect 383514 672618 383546 673174
rect 384102 672618 384134 673174
rect 383514 637174 384134 672618
rect 383514 636618 383546 637174
rect 384102 636618 384134 637174
rect 383514 601174 384134 636618
rect 383514 600618 383546 601174
rect 384102 600618 384134 601174
rect 383514 565174 384134 600618
rect 383514 564618 383546 565174
rect 384102 564618 384134 565174
rect 383514 529174 384134 564618
rect 383514 528618 383546 529174
rect 384102 528618 384134 529174
rect 383514 493174 384134 528618
rect 383514 492618 383546 493174
rect 384102 492618 384134 493174
rect 383514 489603 384134 492618
rect 387234 676894 387854 709082
rect 387234 676338 387266 676894
rect 387822 676338 387854 676894
rect 387234 640894 387854 676338
rect 387234 640338 387266 640894
rect 387822 640338 387854 640894
rect 387234 604894 387854 640338
rect 387234 604338 387266 604894
rect 387822 604338 387854 604894
rect 387234 568894 387854 604338
rect 387234 568338 387266 568894
rect 387822 568338 387854 568894
rect 387234 532894 387854 568338
rect 387234 532338 387266 532894
rect 387822 532338 387854 532894
rect 387234 496894 387854 532338
rect 387234 496338 387266 496894
rect 387822 496338 387854 496894
rect 228954 482058 228986 482614
rect 229542 482058 229574 482614
rect 228954 446614 229574 482058
rect 239208 471454 239528 471486
rect 239208 471218 239250 471454
rect 239486 471218 239528 471454
rect 239208 471134 239528 471218
rect 239208 470898 239250 471134
rect 239486 470898 239528 471134
rect 239208 470866 239528 470898
rect 269928 471454 270248 471486
rect 269928 471218 269970 471454
rect 270206 471218 270248 471454
rect 269928 471134 270248 471218
rect 269928 470898 269970 471134
rect 270206 470898 270248 471134
rect 269928 470866 270248 470898
rect 300648 471454 300968 471486
rect 300648 471218 300690 471454
rect 300926 471218 300968 471454
rect 300648 471134 300968 471218
rect 300648 470898 300690 471134
rect 300926 470898 300968 471134
rect 300648 470866 300968 470898
rect 331368 471454 331688 471486
rect 331368 471218 331410 471454
rect 331646 471218 331688 471454
rect 331368 471134 331688 471218
rect 331368 470898 331410 471134
rect 331646 470898 331688 471134
rect 331368 470866 331688 470898
rect 362088 471454 362408 471486
rect 362088 471218 362130 471454
rect 362366 471218 362408 471454
rect 362088 471134 362408 471218
rect 362088 470898 362130 471134
rect 362366 470898 362408 471134
rect 362088 470866 362408 470898
rect 387234 460894 387854 496338
rect 387234 460338 387266 460894
rect 387822 460338 387854 460894
rect 254568 453454 254888 453486
rect 254568 453218 254610 453454
rect 254846 453218 254888 453454
rect 254568 453134 254888 453218
rect 254568 452898 254610 453134
rect 254846 452898 254888 453134
rect 254568 452866 254888 452898
rect 285288 453454 285608 453486
rect 285288 453218 285330 453454
rect 285566 453218 285608 453454
rect 285288 453134 285608 453218
rect 285288 452898 285330 453134
rect 285566 452898 285608 453134
rect 285288 452866 285608 452898
rect 316008 453454 316328 453486
rect 316008 453218 316050 453454
rect 316286 453218 316328 453454
rect 316008 453134 316328 453218
rect 316008 452898 316050 453134
rect 316286 452898 316328 453134
rect 316008 452866 316328 452898
rect 346728 453454 347048 453486
rect 346728 453218 346770 453454
rect 347006 453218 347048 453454
rect 346728 453134 347048 453218
rect 346728 452898 346770 453134
rect 347006 452898 347048 453134
rect 346728 452866 347048 452898
rect 377448 453454 377768 453486
rect 377448 453218 377490 453454
rect 377726 453218 377768 453454
rect 377448 453134 377768 453218
rect 377448 452898 377490 453134
rect 377726 452898 377768 453134
rect 377448 452866 377768 452898
rect 228954 446058 228986 446614
rect 229542 446058 229574 446614
rect 228954 410614 229574 446058
rect 239208 435454 239528 435486
rect 239208 435218 239250 435454
rect 239486 435218 239528 435454
rect 239208 435134 239528 435218
rect 239208 434898 239250 435134
rect 239486 434898 239528 435134
rect 239208 434866 239528 434898
rect 269928 435454 270248 435486
rect 269928 435218 269970 435454
rect 270206 435218 270248 435454
rect 269928 435134 270248 435218
rect 269928 434898 269970 435134
rect 270206 434898 270248 435134
rect 269928 434866 270248 434898
rect 300648 435454 300968 435486
rect 300648 435218 300690 435454
rect 300926 435218 300968 435454
rect 300648 435134 300968 435218
rect 300648 434898 300690 435134
rect 300926 434898 300968 435134
rect 300648 434866 300968 434898
rect 331368 435454 331688 435486
rect 331368 435218 331410 435454
rect 331646 435218 331688 435454
rect 331368 435134 331688 435218
rect 331368 434898 331410 435134
rect 331646 434898 331688 435134
rect 331368 434866 331688 434898
rect 362088 435454 362408 435486
rect 362088 435218 362130 435454
rect 362366 435218 362408 435454
rect 362088 435134 362408 435218
rect 362088 434898 362130 435134
rect 362366 434898 362408 435134
rect 362088 434866 362408 434898
rect 387234 424894 387854 460338
rect 387234 424338 387266 424894
rect 387822 424338 387854 424894
rect 254568 417454 254888 417486
rect 254568 417218 254610 417454
rect 254846 417218 254888 417454
rect 254568 417134 254888 417218
rect 254568 416898 254610 417134
rect 254846 416898 254888 417134
rect 254568 416866 254888 416898
rect 285288 417454 285608 417486
rect 285288 417218 285330 417454
rect 285566 417218 285608 417454
rect 285288 417134 285608 417218
rect 285288 416898 285330 417134
rect 285566 416898 285608 417134
rect 285288 416866 285608 416898
rect 316008 417454 316328 417486
rect 316008 417218 316050 417454
rect 316286 417218 316328 417454
rect 316008 417134 316328 417218
rect 316008 416898 316050 417134
rect 316286 416898 316328 417134
rect 316008 416866 316328 416898
rect 346728 417454 347048 417486
rect 346728 417218 346770 417454
rect 347006 417218 347048 417454
rect 346728 417134 347048 417218
rect 346728 416898 346770 417134
rect 347006 416898 347048 417134
rect 346728 416866 347048 416898
rect 377448 417454 377768 417486
rect 377448 417218 377490 417454
rect 377726 417218 377768 417454
rect 377448 417134 377768 417218
rect 377448 416898 377490 417134
rect 377726 416898 377768 417134
rect 377448 416866 377768 416898
rect 228954 410058 228986 410614
rect 229542 410058 229574 410614
rect 228954 374614 229574 410058
rect 239208 399454 239528 399486
rect 239208 399218 239250 399454
rect 239486 399218 239528 399454
rect 239208 399134 239528 399218
rect 239208 398898 239250 399134
rect 239486 398898 239528 399134
rect 239208 398866 239528 398898
rect 269928 399454 270248 399486
rect 269928 399218 269970 399454
rect 270206 399218 270248 399454
rect 269928 399134 270248 399218
rect 269928 398898 269970 399134
rect 270206 398898 270248 399134
rect 269928 398866 270248 398898
rect 300648 399454 300968 399486
rect 300648 399218 300690 399454
rect 300926 399218 300968 399454
rect 300648 399134 300968 399218
rect 300648 398898 300690 399134
rect 300926 398898 300968 399134
rect 300648 398866 300968 398898
rect 331368 399454 331688 399486
rect 331368 399218 331410 399454
rect 331646 399218 331688 399454
rect 331368 399134 331688 399218
rect 331368 398898 331410 399134
rect 331646 398898 331688 399134
rect 331368 398866 331688 398898
rect 362088 399454 362408 399486
rect 362088 399218 362130 399454
rect 362366 399218 362408 399454
rect 362088 399134 362408 399218
rect 362088 398898 362130 399134
rect 362366 398898 362408 399134
rect 362088 398866 362408 398898
rect 387234 388894 387854 424338
rect 387234 388338 387266 388894
rect 387822 388338 387854 388894
rect 254568 381454 254888 381486
rect 254568 381218 254610 381454
rect 254846 381218 254888 381454
rect 254568 381134 254888 381218
rect 254568 380898 254610 381134
rect 254846 380898 254888 381134
rect 254568 380866 254888 380898
rect 285288 381454 285608 381486
rect 285288 381218 285330 381454
rect 285566 381218 285608 381454
rect 285288 381134 285608 381218
rect 285288 380898 285330 381134
rect 285566 380898 285608 381134
rect 285288 380866 285608 380898
rect 316008 381454 316328 381486
rect 316008 381218 316050 381454
rect 316286 381218 316328 381454
rect 316008 381134 316328 381218
rect 316008 380898 316050 381134
rect 316286 380898 316328 381134
rect 316008 380866 316328 380898
rect 346728 381454 347048 381486
rect 346728 381218 346770 381454
rect 347006 381218 347048 381454
rect 346728 381134 347048 381218
rect 346728 380898 346770 381134
rect 347006 380898 347048 381134
rect 346728 380866 347048 380898
rect 377448 381454 377768 381486
rect 377448 381218 377490 381454
rect 377726 381218 377768 381454
rect 377448 381134 377768 381218
rect 377448 380898 377490 381134
rect 377726 380898 377768 381134
rect 377448 380866 377768 380898
rect 228954 374058 228986 374614
rect 229542 374058 229574 374614
rect 228954 338614 229574 374058
rect 239208 363454 239528 363486
rect 239208 363218 239250 363454
rect 239486 363218 239528 363454
rect 239208 363134 239528 363218
rect 239208 362898 239250 363134
rect 239486 362898 239528 363134
rect 239208 362866 239528 362898
rect 269928 363454 270248 363486
rect 269928 363218 269970 363454
rect 270206 363218 270248 363454
rect 269928 363134 270248 363218
rect 269928 362898 269970 363134
rect 270206 362898 270248 363134
rect 269928 362866 270248 362898
rect 300648 363454 300968 363486
rect 300648 363218 300690 363454
rect 300926 363218 300968 363454
rect 300648 363134 300968 363218
rect 300648 362898 300690 363134
rect 300926 362898 300968 363134
rect 300648 362866 300968 362898
rect 331368 363454 331688 363486
rect 331368 363218 331410 363454
rect 331646 363218 331688 363454
rect 331368 363134 331688 363218
rect 331368 362898 331410 363134
rect 331646 362898 331688 363134
rect 331368 362866 331688 362898
rect 362088 363454 362408 363486
rect 362088 363218 362130 363454
rect 362366 363218 362408 363454
rect 362088 363134 362408 363218
rect 362088 362898 362130 363134
rect 362366 362898 362408 363134
rect 362088 362866 362408 362898
rect 387234 352894 387854 388338
rect 387234 352338 387266 352894
rect 387822 352338 387854 352894
rect 254568 345454 254888 345486
rect 254568 345218 254610 345454
rect 254846 345218 254888 345454
rect 254568 345134 254888 345218
rect 254568 344898 254610 345134
rect 254846 344898 254888 345134
rect 254568 344866 254888 344898
rect 285288 345454 285608 345486
rect 285288 345218 285330 345454
rect 285566 345218 285608 345454
rect 285288 345134 285608 345218
rect 285288 344898 285330 345134
rect 285566 344898 285608 345134
rect 285288 344866 285608 344898
rect 316008 345454 316328 345486
rect 316008 345218 316050 345454
rect 316286 345218 316328 345454
rect 316008 345134 316328 345218
rect 316008 344898 316050 345134
rect 316286 344898 316328 345134
rect 316008 344866 316328 344898
rect 346728 345454 347048 345486
rect 346728 345218 346770 345454
rect 347006 345218 347048 345454
rect 346728 345134 347048 345218
rect 346728 344898 346770 345134
rect 347006 344898 347048 345134
rect 346728 344866 347048 344898
rect 377448 345454 377768 345486
rect 377448 345218 377490 345454
rect 377726 345218 377768 345454
rect 377448 345134 377768 345218
rect 377448 344898 377490 345134
rect 377726 344898 377768 345134
rect 377448 344866 377768 344898
rect 228954 338058 228986 338614
rect 229542 338058 229574 338614
rect 228954 302614 229574 338058
rect 228954 302058 228986 302614
rect 229542 302058 229574 302614
rect 228954 266614 229574 302058
rect 228954 266058 228986 266614
rect 229542 266058 229574 266614
rect 228954 230614 229574 266058
rect 228954 230058 228986 230614
rect 229542 230058 229574 230614
rect 228954 194614 229574 230058
rect 228954 194058 228986 194614
rect 229542 194058 229574 194614
rect 228954 158614 229574 194058
rect 228954 158058 228986 158614
rect 229542 158058 229574 158614
rect 228954 122614 229574 158058
rect 228954 122058 228986 122614
rect 229542 122058 229574 122614
rect 228954 86614 229574 122058
rect 228954 86058 228986 86614
rect 229542 86058 229574 86614
rect 228954 50614 229574 86058
rect 228954 50058 228986 50614
rect 229542 50058 229574 50614
rect 228954 14614 229574 50058
rect 228954 14058 228986 14614
rect 229542 14058 229574 14614
rect 210954 -7622 210986 -7066
rect 211542 -7622 211574 -7066
rect 210954 -7654 211574 -7622
rect 228954 -6106 229574 14058
rect 235794 309454 236414 336000
rect 235794 308898 235826 309454
rect 236382 308898 236414 309454
rect 235794 273454 236414 308898
rect 235794 272898 235826 273454
rect 236382 272898 236414 273454
rect 235794 237454 236414 272898
rect 235794 236898 235826 237454
rect 236382 236898 236414 237454
rect 235794 201454 236414 236898
rect 235794 200898 235826 201454
rect 236382 200898 236414 201454
rect 235794 165454 236414 200898
rect 235794 164898 235826 165454
rect 236382 164898 236414 165454
rect 235794 129454 236414 164898
rect 235794 128898 235826 129454
rect 236382 128898 236414 129454
rect 235794 93454 236414 128898
rect 235794 92898 235826 93454
rect 236382 92898 236414 93454
rect 235794 57454 236414 92898
rect 235794 56898 235826 57454
rect 236382 56898 236414 57454
rect 235794 21454 236414 56898
rect 235794 20898 235826 21454
rect 236382 20898 236414 21454
rect 235794 -1306 236414 20898
rect 235794 -1862 235826 -1306
rect 236382 -1862 236414 -1306
rect 235794 -1894 236414 -1862
rect 239514 313174 240134 336000
rect 239514 312618 239546 313174
rect 240102 312618 240134 313174
rect 239514 277174 240134 312618
rect 239514 276618 239546 277174
rect 240102 276618 240134 277174
rect 239514 241174 240134 276618
rect 239514 240618 239546 241174
rect 240102 240618 240134 241174
rect 239514 205174 240134 240618
rect 239514 204618 239546 205174
rect 240102 204618 240134 205174
rect 239514 169174 240134 204618
rect 239514 168618 239546 169174
rect 240102 168618 240134 169174
rect 239514 133174 240134 168618
rect 239514 132618 239546 133174
rect 240102 132618 240134 133174
rect 239514 97174 240134 132618
rect 239514 96618 239546 97174
rect 240102 96618 240134 97174
rect 239514 61174 240134 96618
rect 239514 60618 239546 61174
rect 240102 60618 240134 61174
rect 239514 25174 240134 60618
rect 239514 24618 239546 25174
rect 240102 24618 240134 25174
rect 239514 -3226 240134 24618
rect 239514 -3782 239546 -3226
rect 240102 -3782 240134 -3226
rect 239514 -3814 240134 -3782
rect 243234 316894 243854 336000
rect 243234 316338 243266 316894
rect 243822 316338 243854 316894
rect 243234 280894 243854 316338
rect 243234 280338 243266 280894
rect 243822 280338 243854 280894
rect 243234 244894 243854 280338
rect 243234 244338 243266 244894
rect 243822 244338 243854 244894
rect 243234 208894 243854 244338
rect 243234 208338 243266 208894
rect 243822 208338 243854 208894
rect 243234 172894 243854 208338
rect 243234 172338 243266 172894
rect 243822 172338 243854 172894
rect 243234 136894 243854 172338
rect 243234 136338 243266 136894
rect 243822 136338 243854 136894
rect 243234 100894 243854 136338
rect 243234 100338 243266 100894
rect 243822 100338 243854 100894
rect 243234 64894 243854 100338
rect 243234 64338 243266 64894
rect 243822 64338 243854 64894
rect 243234 28894 243854 64338
rect 243234 28338 243266 28894
rect 243822 28338 243854 28894
rect 243234 -5146 243854 28338
rect 243234 -5702 243266 -5146
rect 243822 -5702 243854 -5146
rect 243234 -5734 243854 -5702
rect 246954 320614 247574 336000
rect 246954 320058 246986 320614
rect 247542 320058 247574 320614
rect 246954 284614 247574 320058
rect 246954 284058 246986 284614
rect 247542 284058 247574 284614
rect 246954 248614 247574 284058
rect 246954 248058 246986 248614
rect 247542 248058 247574 248614
rect 246954 212614 247574 248058
rect 246954 212058 246986 212614
rect 247542 212058 247574 212614
rect 246954 176614 247574 212058
rect 246954 176058 246986 176614
rect 247542 176058 247574 176614
rect 246954 140614 247574 176058
rect 246954 140058 246986 140614
rect 247542 140058 247574 140614
rect 246954 104614 247574 140058
rect 246954 104058 246986 104614
rect 247542 104058 247574 104614
rect 246954 68614 247574 104058
rect 246954 68058 246986 68614
rect 247542 68058 247574 68614
rect 246954 32614 247574 68058
rect 246954 32058 246986 32614
rect 247542 32058 247574 32614
rect 228954 -6662 228986 -6106
rect 229542 -6662 229574 -6106
rect 228954 -7654 229574 -6662
rect 246954 -7066 247574 32058
rect 253794 327454 254414 336000
rect 253794 326898 253826 327454
rect 254382 326898 254414 327454
rect 253794 291454 254414 326898
rect 253794 290898 253826 291454
rect 254382 290898 254414 291454
rect 253794 255454 254414 290898
rect 253794 254898 253826 255454
rect 254382 254898 254414 255454
rect 253794 219454 254414 254898
rect 253794 218898 253826 219454
rect 254382 218898 254414 219454
rect 253794 183454 254414 218898
rect 253794 182898 253826 183454
rect 254382 182898 254414 183454
rect 253794 147454 254414 182898
rect 253794 146898 253826 147454
rect 254382 146898 254414 147454
rect 253794 111454 254414 146898
rect 253794 110898 253826 111454
rect 254382 110898 254414 111454
rect 253794 75454 254414 110898
rect 253794 74898 253826 75454
rect 254382 74898 254414 75454
rect 253794 39454 254414 74898
rect 253794 38898 253826 39454
rect 254382 38898 254414 39454
rect 253794 3454 254414 38898
rect 253794 2898 253826 3454
rect 254382 2898 254414 3454
rect 253794 -346 254414 2898
rect 253794 -902 253826 -346
rect 254382 -902 254414 -346
rect 253794 -1894 254414 -902
rect 257514 331174 258134 336000
rect 257514 330618 257546 331174
rect 258102 330618 258134 331174
rect 257514 295174 258134 330618
rect 257514 294618 257546 295174
rect 258102 294618 258134 295174
rect 257514 259174 258134 294618
rect 257514 258618 257546 259174
rect 258102 258618 258134 259174
rect 257514 223174 258134 258618
rect 257514 222618 257546 223174
rect 258102 222618 258134 223174
rect 257514 187174 258134 222618
rect 257514 186618 257546 187174
rect 258102 186618 258134 187174
rect 257514 151174 258134 186618
rect 257514 150618 257546 151174
rect 258102 150618 258134 151174
rect 257514 115174 258134 150618
rect 257514 114618 257546 115174
rect 258102 114618 258134 115174
rect 257514 79174 258134 114618
rect 257514 78618 257546 79174
rect 258102 78618 258134 79174
rect 257514 43174 258134 78618
rect 257514 42618 257546 43174
rect 258102 42618 258134 43174
rect 257514 7174 258134 42618
rect 257514 6618 257546 7174
rect 258102 6618 258134 7174
rect 257514 -2266 258134 6618
rect 257514 -2822 257546 -2266
rect 258102 -2822 258134 -2266
rect 257514 -3814 258134 -2822
rect 261234 334894 261854 336000
rect 261234 334338 261266 334894
rect 261822 334338 261854 334894
rect 261234 298894 261854 334338
rect 261234 298338 261266 298894
rect 261822 298338 261854 298894
rect 261234 262894 261854 298338
rect 261234 262338 261266 262894
rect 261822 262338 261854 262894
rect 261234 226894 261854 262338
rect 261234 226338 261266 226894
rect 261822 226338 261854 226894
rect 261234 190894 261854 226338
rect 261234 190338 261266 190894
rect 261822 190338 261854 190894
rect 261234 154894 261854 190338
rect 261234 154338 261266 154894
rect 261822 154338 261854 154894
rect 261234 118894 261854 154338
rect 261234 118338 261266 118894
rect 261822 118338 261854 118894
rect 261234 82894 261854 118338
rect 261234 82338 261266 82894
rect 261822 82338 261854 82894
rect 261234 46894 261854 82338
rect 261234 46338 261266 46894
rect 261822 46338 261854 46894
rect 261234 10894 261854 46338
rect 261234 10338 261266 10894
rect 261822 10338 261854 10894
rect 261234 -4186 261854 10338
rect 261234 -4742 261266 -4186
rect 261822 -4742 261854 -4186
rect 261234 -5734 261854 -4742
rect 264954 302614 265574 336000
rect 264954 302058 264986 302614
rect 265542 302058 265574 302614
rect 264954 266614 265574 302058
rect 264954 266058 264986 266614
rect 265542 266058 265574 266614
rect 264954 230614 265574 266058
rect 264954 230058 264986 230614
rect 265542 230058 265574 230614
rect 264954 194614 265574 230058
rect 264954 194058 264986 194614
rect 265542 194058 265574 194614
rect 264954 158614 265574 194058
rect 264954 158058 264986 158614
rect 265542 158058 265574 158614
rect 264954 122614 265574 158058
rect 264954 122058 264986 122614
rect 265542 122058 265574 122614
rect 264954 86614 265574 122058
rect 264954 86058 264986 86614
rect 265542 86058 265574 86614
rect 264954 50614 265574 86058
rect 264954 50058 264986 50614
rect 265542 50058 265574 50614
rect 264954 14614 265574 50058
rect 264954 14058 264986 14614
rect 265542 14058 265574 14614
rect 246954 -7622 246986 -7066
rect 247542 -7622 247574 -7066
rect 246954 -7654 247574 -7622
rect 264954 -6106 265574 14058
rect 271794 309454 272414 336000
rect 271794 308898 271826 309454
rect 272382 308898 272414 309454
rect 271794 273454 272414 308898
rect 271794 272898 271826 273454
rect 272382 272898 272414 273454
rect 271794 237454 272414 272898
rect 271794 236898 271826 237454
rect 272382 236898 272414 237454
rect 271794 201454 272414 236898
rect 271794 200898 271826 201454
rect 272382 200898 272414 201454
rect 271794 165454 272414 200898
rect 271794 164898 271826 165454
rect 272382 164898 272414 165454
rect 271794 129454 272414 164898
rect 271794 128898 271826 129454
rect 272382 128898 272414 129454
rect 271794 93454 272414 128898
rect 271794 92898 271826 93454
rect 272382 92898 272414 93454
rect 271794 57454 272414 92898
rect 271794 56898 271826 57454
rect 272382 56898 272414 57454
rect 271794 21454 272414 56898
rect 271794 20898 271826 21454
rect 272382 20898 272414 21454
rect 271794 -1306 272414 20898
rect 271794 -1862 271826 -1306
rect 272382 -1862 272414 -1306
rect 271794 -1894 272414 -1862
rect 275514 313174 276134 336000
rect 275514 312618 275546 313174
rect 276102 312618 276134 313174
rect 275514 277174 276134 312618
rect 275514 276618 275546 277174
rect 276102 276618 276134 277174
rect 275514 241174 276134 276618
rect 275514 240618 275546 241174
rect 276102 240618 276134 241174
rect 275514 205174 276134 240618
rect 275514 204618 275546 205174
rect 276102 204618 276134 205174
rect 275514 169174 276134 204618
rect 275514 168618 275546 169174
rect 276102 168618 276134 169174
rect 275514 133174 276134 168618
rect 275514 132618 275546 133174
rect 276102 132618 276134 133174
rect 275514 97174 276134 132618
rect 275514 96618 275546 97174
rect 276102 96618 276134 97174
rect 275514 61174 276134 96618
rect 275514 60618 275546 61174
rect 276102 60618 276134 61174
rect 275514 25174 276134 60618
rect 275514 24618 275546 25174
rect 276102 24618 276134 25174
rect 275514 -3226 276134 24618
rect 275514 -3782 275546 -3226
rect 276102 -3782 276134 -3226
rect 275514 -3814 276134 -3782
rect 279234 316894 279854 336000
rect 279234 316338 279266 316894
rect 279822 316338 279854 316894
rect 279234 280894 279854 316338
rect 279234 280338 279266 280894
rect 279822 280338 279854 280894
rect 279234 244894 279854 280338
rect 279234 244338 279266 244894
rect 279822 244338 279854 244894
rect 279234 208894 279854 244338
rect 279234 208338 279266 208894
rect 279822 208338 279854 208894
rect 279234 172894 279854 208338
rect 279234 172338 279266 172894
rect 279822 172338 279854 172894
rect 279234 136894 279854 172338
rect 279234 136338 279266 136894
rect 279822 136338 279854 136894
rect 279234 100894 279854 136338
rect 279234 100338 279266 100894
rect 279822 100338 279854 100894
rect 279234 64894 279854 100338
rect 279234 64338 279266 64894
rect 279822 64338 279854 64894
rect 279234 28894 279854 64338
rect 279234 28338 279266 28894
rect 279822 28338 279854 28894
rect 279234 -5146 279854 28338
rect 279234 -5702 279266 -5146
rect 279822 -5702 279854 -5146
rect 279234 -5734 279854 -5702
rect 282954 320614 283574 336000
rect 282954 320058 282986 320614
rect 283542 320058 283574 320614
rect 282954 284614 283574 320058
rect 282954 284058 282986 284614
rect 283542 284058 283574 284614
rect 282954 248614 283574 284058
rect 282954 248058 282986 248614
rect 283542 248058 283574 248614
rect 282954 212614 283574 248058
rect 282954 212058 282986 212614
rect 283542 212058 283574 212614
rect 282954 176614 283574 212058
rect 282954 176058 282986 176614
rect 283542 176058 283574 176614
rect 282954 140614 283574 176058
rect 282954 140058 282986 140614
rect 283542 140058 283574 140614
rect 282954 104614 283574 140058
rect 282954 104058 282986 104614
rect 283542 104058 283574 104614
rect 282954 68614 283574 104058
rect 282954 68058 282986 68614
rect 283542 68058 283574 68614
rect 282954 32614 283574 68058
rect 282954 32058 282986 32614
rect 283542 32058 283574 32614
rect 264954 -6662 264986 -6106
rect 265542 -6662 265574 -6106
rect 264954 -7654 265574 -6662
rect 282954 -7066 283574 32058
rect 289794 327454 290414 336000
rect 289794 326898 289826 327454
rect 290382 326898 290414 327454
rect 289794 291454 290414 326898
rect 289794 290898 289826 291454
rect 290382 290898 290414 291454
rect 289794 255454 290414 290898
rect 289794 254898 289826 255454
rect 290382 254898 290414 255454
rect 289794 219454 290414 254898
rect 289794 218898 289826 219454
rect 290382 218898 290414 219454
rect 289794 183454 290414 218898
rect 289794 182898 289826 183454
rect 290382 182898 290414 183454
rect 289794 147454 290414 182898
rect 289794 146898 289826 147454
rect 290382 146898 290414 147454
rect 289794 111454 290414 146898
rect 289794 110898 289826 111454
rect 290382 110898 290414 111454
rect 289794 75454 290414 110898
rect 289794 74898 289826 75454
rect 290382 74898 290414 75454
rect 289794 39454 290414 74898
rect 289794 38898 289826 39454
rect 290382 38898 290414 39454
rect 289794 3454 290414 38898
rect 289794 2898 289826 3454
rect 290382 2898 290414 3454
rect 289794 -346 290414 2898
rect 289794 -902 289826 -346
rect 290382 -902 290414 -346
rect 289794 -1894 290414 -902
rect 293514 331174 294134 336000
rect 293514 330618 293546 331174
rect 294102 330618 294134 331174
rect 293514 295174 294134 330618
rect 293514 294618 293546 295174
rect 294102 294618 294134 295174
rect 293514 259174 294134 294618
rect 293514 258618 293546 259174
rect 294102 258618 294134 259174
rect 293514 223174 294134 258618
rect 293514 222618 293546 223174
rect 294102 222618 294134 223174
rect 293514 187174 294134 222618
rect 293514 186618 293546 187174
rect 294102 186618 294134 187174
rect 293514 151174 294134 186618
rect 293514 150618 293546 151174
rect 294102 150618 294134 151174
rect 293514 115174 294134 150618
rect 293514 114618 293546 115174
rect 294102 114618 294134 115174
rect 293514 79174 294134 114618
rect 293514 78618 293546 79174
rect 294102 78618 294134 79174
rect 293514 43174 294134 78618
rect 293514 42618 293546 43174
rect 294102 42618 294134 43174
rect 293514 7174 294134 42618
rect 293514 6618 293546 7174
rect 294102 6618 294134 7174
rect 293514 -2266 294134 6618
rect 293514 -2822 293546 -2266
rect 294102 -2822 294134 -2266
rect 293514 -3814 294134 -2822
rect 297234 334894 297854 336000
rect 297234 334338 297266 334894
rect 297822 334338 297854 334894
rect 297234 298894 297854 334338
rect 297234 298338 297266 298894
rect 297822 298338 297854 298894
rect 297234 262894 297854 298338
rect 297234 262338 297266 262894
rect 297822 262338 297854 262894
rect 297234 226894 297854 262338
rect 297234 226338 297266 226894
rect 297822 226338 297854 226894
rect 297234 190894 297854 226338
rect 297234 190338 297266 190894
rect 297822 190338 297854 190894
rect 297234 154894 297854 190338
rect 297234 154338 297266 154894
rect 297822 154338 297854 154894
rect 297234 118894 297854 154338
rect 297234 118338 297266 118894
rect 297822 118338 297854 118894
rect 297234 82894 297854 118338
rect 297234 82338 297266 82894
rect 297822 82338 297854 82894
rect 297234 46894 297854 82338
rect 297234 46338 297266 46894
rect 297822 46338 297854 46894
rect 297234 10894 297854 46338
rect 297234 10338 297266 10894
rect 297822 10338 297854 10894
rect 297234 -4186 297854 10338
rect 297234 -4742 297266 -4186
rect 297822 -4742 297854 -4186
rect 297234 -5734 297854 -4742
rect 300954 302614 301574 336000
rect 300954 302058 300986 302614
rect 301542 302058 301574 302614
rect 300954 266614 301574 302058
rect 300954 266058 300986 266614
rect 301542 266058 301574 266614
rect 300954 230614 301574 266058
rect 300954 230058 300986 230614
rect 301542 230058 301574 230614
rect 300954 194614 301574 230058
rect 300954 194058 300986 194614
rect 301542 194058 301574 194614
rect 300954 158614 301574 194058
rect 300954 158058 300986 158614
rect 301542 158058 301574 158614
rect 300954 122614 301574 158058
rect 300954 122058 300986 122614
rect 301542 122058 301574 122614
rect 300954 86614 301574 122058
rect 300954 86058 300986 86614
rect 301542 86058 301574 86614
rect 300954 50614 301574 86058
rect 300954 50058 300986 50614
rect 301542 50058 301574 50614
rect 300954 14614 301574 50058
rect 300954 14058 300986 14614
rect 301542 14058 301574 14614
rect 282954 -7622 282986 -7066
rect 283542 -7622 283574 -7066
rect 282954 -7654 283574 -7622
rect 300954 -6106 301574 14058
rect 307794 309454 308414 336000
rect 307794 308898 307826 309454
rect 308382 308898 308414 309454
rect 307794 273454 308414 308898
rect 307794 272898 307826 273454
rect 308382 272898 308414 273454
rect 307794 237454 308414 272898
rect 307794 236898 307826 237454
rect 308382 236898 308414 237454
rect 307794 201454 308414 236898
rect 307794 200898 307826 201454
rect 308382 200898 308414 201454
rect 307794 165454 308414 200898
rect 307794 164898 307826 165454
rect 308382 164898 308414 165454
rect 307794 129454 308414 164898
rect 307794 128898 307826 129454
rect 308382 128898 308414 129454
rect 307794 93454 308414 128898
rect 307794 92898 307826 93454
rect 308382 92898 308414 93454
rect 307794 57454 308414 92898
rect 307794 56898 307826 57454
rect 308382 56898 308414 57454
rect 307794 21454 308414 56898
rect 307794 20898 307826 21454
rect 308382 20898 308414 21454
rect 307794 -1306 308414 20898
rect 307794 -1862 307826 -1306
rect 308382 -1862 308414 -1306
rect 307794 -1894 308414 -1862
rect 311514 313174 312134 336000
rect 311514 312618 311546 313174
rect 312102 312618 312134 313174
rect 311514 277174 312134 312618
rect 311514 276618 311546 277174
rect 312102 276618 312134 277174
rect 311514 241174 312134 276618
rect 311514 240618 311546 241174
rect 312102 240618 312134 241174
rect 311514 205174 312134 240618
rect 311514 204618 311546 205174
rect 312102 204618 312134 205174
rect 311514 169174 312134 204618
rect 311514 168618 311546 169174
rect 312102 168618 312134 169174
rect 311514 133174 312134 168618
rect 311514 132618 311546 133174
rect 312102 132618 312134 133174
rect 311514 97174 312134 132618
rect 311514 96618 311546 97174
rect 312102 96618 312134 97174
rect 311514 61174 312134 96618
rect 311514 60618 311546 61174
rect 312102 60618 312134 61174
rect 311514 25174 312134 60618
rect 311514 24618 311546 25174
rect 312102 24618 312134 25174
rect 311514 -3226 312134 24618
rect 311514 -3782 311546 -3226
rect 312102 -3782 312134 -3226
rect 311514 -3814 312134 -3782
rect 315234 316894 315854 336000
rect 315234 316338 315266 316894
rect 315822 316338 315854 316894
rect 315234 280894 315854 316338
rect 315234 280338 315266 280894
rect 315822 280338 315854 280894
rect 315234 244894 315854 280338
rect 315234 244338 315266 244894
rect 315822 244338 315854 244894
rect 315234 208894 315854 244338
rect 315234 208338 315266 208894
rect 315822 208338 315854 208894
rect 315234 172894 315854 208338
rect 315234 172338 315266 172894
rect 315822 172338 315854 172894
rect 315234 136894 315854 172338
rect 315234 136338 315266 136894
rect 315822 136338 315854 136894
rect 315234 100894 315854 136338
rect 315234 100338 315266 100894
rect 315822 100338 315854 100894
rect 315234 64894 315854 100338
rect 315234 64338 315266 64894
rect 315822 64338 315854 64894
rect 315234 28894 315854 64338
rect 315234 28338 315266 28894
rect 315822 28338 315854 28894
rect 315234 -5146 315854 28338
rect 315234 -5702 315266 -5146
rect 315822 -5702 315854 -5146
rect 315234 -5734 315854 -5702
rect 318954 320614 319574 336000
rect 318954 320058 318986 320614
rect 319542 320058 319574 320614
rect 318954 284614 319574 320058
rect 318954 284058 318986 284614
rect 319542 284058 319574 284614
rect 318954 248614 319574 284058
rect 318954 248058 318986 248614
rect 319542 248058 319574 248614
rect 318954 212614 319574 248058
rect 318954 212058 318986 212614
rect 319542 212058 319574 212614
rect 318954 176614 319574 212058
rect 318954 176058 318986 176614
rect 319542 176058 319574 176614
rect 318954 140614 319574 176058
rect 318954 140058 318986 140614
rect 319542 140058 319574 140614
rect 318954 104614 319574 140058
rect 318954 104058 318986 104614
rect 319542 104058 319574 104614
rect 318954 68614 319574 104058
rect 318954 68058 318986 68614
rect 319542 68058 319574 68614
rect 318954 32614 319574 68058
rect 318954 32058 318986 32614
rect 319542 32058 319574 32614
rect 300954 -6662 300986 -6106
rect 301542 -6662 301574 -6106
rect 300954 -7654 301574 -6662
rect 318954 -7066 319574 32058
rect 325794 327454 326414 336000
rect 325794 326898 325826 327454
rect 326382 326898 326414 327454
rect 325794 291454 326414 326898
rect 325794 290898 325826 291454
rect 326382 290898 326414 291454
rect 325794 255454 326414 290898
rect 325794 254898 325826 255454
rect 326382 254898 326414 255454
rect 325794 219454 326414 254898
rect 325794 218898 325826 219454
rect 326382 218898 326414 219454
rect 325794 183454 326414 218898
rect 325794 182898 325826 183454
rect 326382 182898 326414 183454
rect 325794 147454 326414 182898
rect 325794 146898 325826 147454
rect 326382 146898 326414 147454
rect 325794 111454 326414 146898
rect 325794 110898 325826 111454
rect 326382 110898 326414 111454
rect 325794 75454 326414 110898
rect 325794 74898 325826 75454
rect 326382 74898 326414 75454
rect 325794 39454 326414 74898
rect 325794 38898 325826 39454
rect 326382 38898 326414 39454
rect 325794 3454 326414 38898
rect 325794 2898 325826 3454
rect 326382 2898 326414 3454
rect 325794 -346 326414 2898
rect 325794 -902 325826 -346
rect 326382 -902 326414 -346
rect 325794 -1894 326414 -902
rect 329514 331174 330134 336000
rect 329514 330618 329546 331174
rect 330102 330618 330134 331174
rect 329514 295174 330134 330618
rect 329514 294618 329546 295174
rect 330102 294618 330134 295174
rect 329514 259174 330134 294618
rect 329514 258618 329546 259174
rect 330102 258618 330134 259174
rect 329514 223174 330134 258618
rect 329514 222618 329546 223174
rect 330102 222618 330134 223174
rect 329514 187174 330134 222618
rect 329514 186618 329546 187174
rect 330102 186618 330134 187174
rect 329514 151174 330134 186618
rect 329514 150618 329546 151174
rect 330102 150618 330134 151174
rect 329514 115174 330134 150618
rect 329514 114618 329546 115174
rect 330102 114618 330134 115174
rect 329514 79174 330134 114618
rect 329514 78618 329546 79174
rect 330102 78618 330134 79174
rect 329514 43174 330134 78618
rect 329514 42618 329546 43174
rect 330102 42618 330134 43174
rect 329514 7174 330134 42618
rect 329514 6618 329546 7174
rect 330102 6618 330134 7174
rect 329514 -2266 330134 6618
rect 329514 -2822 329546 -2266
rect 330102 -2822 330134 -2266
rect 329514 -3814 330134 -2822
rect 333234 334894 333854 336000
rect 333234 334338 333266 334894
rect 333822 334338 333854 334894
rect 333234 298894 333854 334338
rect 333234 298338 333266 298894
rect 333822 298338 333854 298894
rect 333234 262894 333854 298338
rect 333234 262338 333266 262894
rect 333822 262338 333854 262894
rect 333234 226894 333854 262338
rect 333234 226338 333266 226894
rect 333822 226338 333854 226894
rect 333234 190894 333854 226338
rect 333234 190338 333266 190894
rect 333822 190338 333854 190894
rect 333234 154894 333854 190338
rect 333234 154338 333266 154894
rect 333822 154338 333854 154894
rect 333234 118894 333854 154338
rect 333234 118338 333266 118894
rect 333822 118338 333854 118894
rect 333234 82894 333854 118338
rect 333234 82338 333266 82894
rect 333822 82338 333854 82894
rect 333234 46894 333854 82338
rect 333234 46338 333266 46894
rect 333822 46338 333854 46894
rect 333234 10894 333854 46338
rect 333234 10338 333266 10894
rect 333822 10338 333854 10894
rect 333234 -4186 333854 10338
rect 333234 -4742 333266 -4186
rect 333822 -4742 333854 -4186
rect 333234 -5734 333854 -4742
rect 336954 302614 337574 336000
rect 336954 302058 336986 302614
rect 337542 302058 337574 302614
rect 336954 266614 337574 302058
rect 336954 266058 336986 266614
rect 337542 266058 337574 266614
rect 336954 230614 337574 266058
rect 336954 230058 336986 230614
rect 337542 230058 337574 230614
rect 336954 194614 337574 230058
rect 336954 194058 336986 194614
rect 337542 194058 337574 194614
rect 336954 158614 337574 194058
rect 336954 158058 336986 158614
rect 337542 158058 337574 158614
rect 336954 122614 337574 158058
rect 336954 122058 336986 122614
rect 337542 122058 337574 122614
rect 336954 86614 337574 122058
rect 336954 86058 336986 86614
rect 337542 86058 337574 86614
rect 336954 50614 337574 86058
rect 336954 50058 336986 50614
rect 337542 50058 337574 50614
rect 336954 14614 337574 50058
rect 336954 14058 336986 14614
rect 337542 14058 337574 14614
rect 318954 -7622 318986 -7066
rect 319542 -7622 319574 -7066
rect 318954 -7654 319574 -7622
rect 336954 -6106 337574 14058
rect 343794 309454 344414 336000
rect 343794 308898 343826 309454
rect 344382 308898 344414 309454
rect 343794 273454 344414 308898
rect 343794 272898 343826 273454
rect 344382 272898 344414 273454
rect 343794 237454 344414 272898
rect 343794 236898 343826 237454
rect 344382 236898 344414 237454
rect 343794 201454 344414 236898
rect 343794 200898 343826 201454
rect 344382 200898 344414 201454
rect 343794 165454 344414 200898
rect 343794 164898 343826 165454
rect 344382 164898 344414 165454
rect 343794 129454 344414 164898
rect 343794 128898 343826 129454
rect 344382 128898 344414 129454
rect 343794 93454 344414 128898
rect 343794 92898 343826 93454
rect 344382 92898 344414 93454
rect 343794 57454 344414 92898
rect 343794 56898 343826 57454
rect 344382 56898 344414 57454
rect 343794 21454 344414 56898
rect 343794 20898 343826 21454
rect 344382 20898 344414 21454
rect 343794 -1306 344414 20898
rect 343794 -1862 343826 -1306
rect 344382 -1862 344414 -1306
rect 343794 -1894 344414 -1862
rect 347514 313174 348134 336000
rect 347514 312618 347546 313174
rect 348102 312618 348134 313174
rect 347514 277174 348134 312618
rect 347514 276618 347546 277174
rect 348102 276618 348134 277174
rect 347514 241174 348134 276618
rect 347514 240618 347546 241174
rect 348102 240618 348134 241174
rect 347514 205174 348134 240618
rect 347514 204618 347546 205174
rect 348102 204618 348134 205174
rect 347514 169174 348134 204618
rect 347514 168618 347546 169174
rect 348102 168618 348134 169174
rect 347514 133174 348134 168618
rect 347514 132618 347546 133174
rect 348102 132618 348134 133174
rect 347514 97174 348134 132618
rect 347514 96618 347546 97174
rect 348102 96618 348134 97174
rect 347514 61174 348134 96618
rect 347514 60618 347546 61174
rect 348102 60618 348134 61174
rect 347514 25174 348134 60618
rect 347514 24618 347546 25174
rect 348102 24618 348134 25174
rect 347514 -3226 348134 24618
rect 347514 -3782 347546 -3226
rect 348102 -3782 348134 -3226
rect 347514 -3814 348134 -3782
rect 351234 316894 351854 336000
rect 351234 316338 351266 316894
rect 351822 316338 351854 316894
rect 351234 280894 351854 316338
rect 351234 280338 351266 280894
rect 351822 280338 351854 280894
rect 351234 244894 351854 280338
rect 351234 244338 351266 244894
rect 351822 244338 351854 244894
rect 351234 208894 351854 244338
rect 351234 208338 351266 208894
rect 351822 208338 351854 208894
rect 351234 172894 351854 208338
rect 351234 172338 351266 172894
rect 351822 172338 351854 172894
rect 351234 136894 351854 172338
rect 351234 136338 351266 136894
rect 351822 136338 351854 136894
rect 351234 100894 351854 136338
rect 351234 100338 351266 100894
rect 351822 100338 351854 100894
rect 351234 64894 351854 100338
rect 351234 64338 351266 64894
rect 351822 64338 351854 64894
rect 351234 28894 351854 64338
rect 351234 28338 351266 28894
rect 351822 28338 351854 28894
rect 351234 -5146 351854 28338
rect 351234 -5702 351266 -5146
rect 351822 -5702 351854 -5146
rect 351234 -5734 351854 -5702
rect 354954 320614 355574 336000
rect 354954 320058 354986 320614
rect 355542 320058 355574 320614
rect 354954 284614 355574 320058
rect 354954 284058 354986 284614
rect 355542 284058 355574 284614
rect 354954 248614 355574 284058
rect 354954 248058 354986 248614
rect 355542 248058 355574 248614
rect 354954 212614 355574 248058
rect 354954 212058 354986 212614
rect 355542 212058 355574 212614
rect 354954 176614 355574 212058
rect 354954 176058 354986 176614
rect 355542 176058 355574 176614
rect 354954 140614 355574 176058
rect 354954 140058 354986 140614
rect 355542 140058 355574 140614
rect 354954 104614 355574 140058
rect 354954 104058 354986 104614
rect 355542 104058 355574 104614
rect 354954 68614 355574 104058
rect 354954 68058 354986 68614
rect 355542 68058 355574 68614
rect 354954 32614 355574 68058
rect 354954 32058 354986 32614
rect 355542 32058 355574 32614
rect 336954 -6662 336986 -6106
rect 337542 -6662 337574 -6106
rect 336954 -7654 337574 -6662
rect 354954 -7066 355574 32058
rect 361794 327454 362414 336000
rect 361794 326898 361826 327454
rect 362382 326898 362414 327454
rect 361794 291454 362414 326898
rect 361794 290898 361826 291454
rect 362382 290898 362414 291454
rect 361794 255454 362414 290898
rect 361794 254898 361826 255454
rect 362382 254898 362414 255454
rect 361794 219454 362414 254898
rect 361794 218898 361826 219454
rect 362382 218898 362414 219454
rect 361794 183454 362414 218898
rect 361794 182898 361826 183454
rect 362382 182898 362414 183454
rect 361794 147454 362414 182898
rect 361794 146898 361826 147454
rect 362382 146898 362414 147454
rect 361794 111454 362414 146898
rect 361794 110898 361826 111454
rect 362382 110898 362414 111454
rect 361794 75454 362414 110898
rect 361794 74898 361826 75454
rect 362382 74898 362414 75454
rect 361794 39454 362414 74898
rect 361794 38898 361826 39454
rect 362382 38898 362414 39454
rect 361794 3454 362414 38898
rect 361794 2898 361826 3454
rect 362382 2898 362414 3454
rect 361794 -346 362414 2898
rect 361794 -902 361826 -346
rect 362382 -902 362414 -346
rect 361794 -1894 362414 -902
rect 365514 331174 366134 336000
rect 365514 330618 365546 331174
rect 366102 330618 366134 331174
rect 365514 295174 366134 330618
rect 365514 294618 365546 295174
rect 366102 294618 366134 295174
rect 365514 259174 366134 294618
rect 365514 258618 365546 259174
rect 366102 258618 366134 259174
rect 365514 223174 366134 258618
rect 365514 222618 365546 223174
rect 366102 222618 366134 223174
rect 365514 187174 366134 222618
rect 365514 186618 365546 187174
rect 366102 186618 366134 187174
rect 365514 151174 366134 186618
rect 365514 150618 365546 151174
rect 366102 150618 366134 151174
rect 365514 115174 366134 150618
rect 365514 114618 365546 115174
rect 366102 114618 366134 115174
rect 365514 79174 366134 114618
rect 365514 78618 365546 79174
rect 366102 78618 366134 79174
rect 365514 43174 366134 78618
rect 365514 42618 365546 43174
rect 366102 42618 366134 43174
rect 365514 7174 366134 42618
rect 365514 6618 365546 7174
rect 366102 6618 366134 7174
rect 365514 -2266 366134 6618
rect 365514 -2822 365546 -2266
rect 366102 -2822 366134 -2266
rect 365514 -3814 366134 -2822
rect 369234 334894 369854 336000
rect 369234 334338 369266 334894
rect 369822 334338 369854 334894
rect 369234 298894 369854 334338
rect 369234 298338 369266 298894
rect 369822 298338 369854 298894
rect 369234 262894 369854 298338
rect 369234 262338 369266 262894
rect 369822 262338 369854 262894
rect 369234 226894 369854 262338
rect 369234 226338 369266 226894
rect 369822 226338 369854 226894
rect 369234 190894 369854 226338
rect 369234 190338 369266 190894
rect 369822 190338 369854 190894
rect 369234 154894 369854 190338
rect 369234 154338 369266 154894
rect 369822 154338 369854 154894
rect 369234 118894 369854 154338
rect 369234 118338 369266 118894
rect 369822 118338 369854 118894
rect 369234 82894 369854 118338
rect 369234 82338 369266 82894
rect 369822 82338 369854 82894
rect 369234 46894 369854 82338
rect 369234 46338 369266 46894
rect 369822 46338 369854 46894
rect 369234 10894 369854 46338
rect 369234 10338 369266 10894
rect 369822 10338 369854 10894
rect 369234 -4186 369854 10338
rect 369234 -4742 369266 -4186
rect 369822 -4742 369854 -4186
rect 369234 -5734 369854 -4742
rect 372954 302614 373574 336000
rect 372954 302058 372986 302614
rect 373542 302058 373574 302614
rect 372954 266614 373574 302058
rect 372954 266058 372986 266614
rect 373542 266058 373574 266614
rect 372954 230614 373574 266058
rect 372954 230058 372986 230614
rect 373542 230058 373574 230614
rect 372954 194614 373574 230058
rect 372954 194058 372986 194614
rect 373542 194058 373574 194614
rect 372954 158614 373574 194058
rect 372954 158058 372986 158614
rect 373542 158058 373574 158614
rect 372954 122614 373574 158058
rect 372954 122058 372986 122614
rect 373542 122058 373574 122614
rect 372954 86614 373574 122058
rect 372954 86058 372986 86614
rect 373542 86058 373574 86614
rect 372954 50614 373574 86058
rect 372954 50058 372986 50614
rect 373542 50058 373574 50614
rect 372954 14614 373574 50058
rect 372954 14058 372986 14614
rect 373542 14058 373574 14614
rect 354954 -7622 354986 -7066
rect 355542 -7622 355574 -7066
rect 354954 -7654 355574 -7622
rect 372954 -6106 373574 14058
rect 379794 309454 380414 336000
rect 379794 308898 379826 309454
rect 380382 308898 380414 309454
rect 379794 273454 380414 308898
rect 379794 272898 379826 273454
rect 380382 272898 380414 273454
rect 379794 237454 380414 272898
rect 379794 236898 379826 237454
rect 380382 236898 380414 237454
rect 379794 201454 380414 236898
rect 379794 200898 379826 201454
rect 380382 200898 380414 201454
rect 379794 165454 380414 200898
rect 379794 164898 379826 165454
rect 380382 164898 380414 165454
rect 379794 129454 380414 164898
rect 379794 128898 379826 129454
rect 380382 128898 380414 129454
rect 379794 93454 380414 128898
rect 379794 92898 379826 93454
rect 380382 92898 380414 93454
rect 379794 57454 380414 92898
rect 379794 56898 379826 57454
rect 380382 56898 380414 57454
rect 379794 21454 380414 56898
rect 379794 20898 379826 21454
rect 380382 20898 380414 21454
rect 379794 -1306 380414 20898
rect 379794 -1862 379826 -1306
rect 380382 -1862 380414 -1306
rect 379794 -1894 380414 -1862
rect 383514 313174 384134 336000
rect 383514 312618 383546 313174
rect 384102 312618 384134 313174
rect 383514 277174 384134 312618
rect 383514 276618 383546 277174
rect 384102 276618 384134 277174
rect 383514 241174 384134 276618
rect 383514 240618 383546 241174
rect 384102 240618 384134 241174
rect 383514 205174 384134 240618
rect 383514 204618 383546 205174
rect 384102 204618 384134 205174
rect 383514 169174 384134 204618
rect 383514 168618 383546 169174
rect 384102 168618 384134 169174
rect 383514 133174 384134 168618
rect 383514 132618 383546 133174
rect 384102 132618 384134 133174
rect 383514 97174 384134 132618
rect 383514 96618 383546 97174
rect 384102 96618 384134 97174
rect 383514 61174 384134 96618
rect 383514 60618 383546 61174
rect 384102 60618 384134 61174
rect 383514 25174 384134 60618
rect 383514 24618 383546 25174
rect 384102 24618 384134 25174
rect 383514 -3226 384134 24618
rect 383514 -3782 383546 -3226
rect 384102 -3782 384134 -3226
rect 383514 -3814 384134 -3782
rect 387234 316894 387854 352338
rect 387234 316338 387266 316894
rect 387822 316338 387854 316894
rect 387234 280894 387854 316338
rect 387234 280338 387266 280894
rect 387822 280338 387854 280894
rect 387234 244894 387854 280338
rect 387234 244338 387266 244894
rect 387822 244338 387854 244894
rect 387234 208894 387854 244338
rect 387234 208338 387266 208894
rect 387822 208338 387854 208894
rect 387234 172894 387854 208338
rect 387234 172338 387266 172894
rect 387822 172338 387854 172894
rect 387234 136894 387854 172338
rect 387234 136338 387266 136894
rect 387822 136338 387854 136894
rect 387234 100894 387854 136338
rect 387234 100338 387266 100894
rect 387822 100338 387854 100894
rect 387234 64894 387854 100338
rect 387234 64338 387266 64894
rect 387822 64338 387854 64894
rect 387234 28894 387854 64338
rect 387234 28338 387266 28894
rect 387822 28338 387854 28894
rect 387234 -5146 387854 28338
rect 387234 -5702 387266 -5146
rect 387822 -5702 387854 -5146
rect 387234 -5734 387854 -5702
rect 390954 680614 391574 711002
rect 408954 710598 409574 711590
rect 408954 710042 408986 710598
rect 409542 710042 409574 710598
rect 405234 708678 405854 709670
rect 405234 708122 405266 708678
rect 405822 708122 405854 708678
rect 401514 706758 402134 707750
rect 401514 706202 401546 706758
rect 402102 706202 402134 706758
rect 390954 680058 390986 680614
rect 391542 680058 391574 680614
rect 390954 644614 391574 680058
rect 390954 644058 390986 644614
rect 391542 644058 391574 644614
rect 390954 608614 391574 644058
rect 390954 608058 390986 608614
rect 391542 608058 391574 608614
rect 390954 572614 391574 608058
rect 390954 572058 390986 572614
rect 391542 572058 391574 572614
rect 390954 536614 391574 572058
rect 390954 536058 390986 536614
rect 391542 536058 391574 536614
rect 390954 500614 391574 536058
rect 390954 500058 390986 500614
rect 391542 500058 391574 500614
rect 390954 464614 391574 500058
rect 390954 464058 390986 464614
rect 391542 464058 391574 464614
rect 390954 428614 391574 464058
rect 390954 428058 390986 428614
rect 391542 428058 391574 428614
rect 390954 392614 391574 428058
rect 390954 392058 390986 392614
rect 391542 392058 391574 392614
rect 390954 356614 391574 392058
rect 390954 356058 390986 356614
rect 391542 356058 391574 356614
rect 390954 320614 391574 356058
rect 390954 320058 390986 320614
rect 391542 320058 391574 320614
rect 390954 284614 391574 320058
rect 390954 284058 390986 284614
rect 391542 284058 391574 284614
rect 390954 248614 391574 284058
rect 390954 248058 390986 248614
rect 391542 248058 391574 248614
rect 390954 212614 391574 248058
rect 390954 212058 390986 212614
rect 391542 212058 391574 212614
rect 390954 176614 391574 212058
rect 390954 176058 390986 176614
rect 391542 176058 391574 176614
rect 390954 140614 391574 176058
rect 390954 140058 390986 140614
rect 391542 140058 391574 140614
rect 390954 104614 391574 140058
rect 390954 104058 390986 104614
rect 391542 104058 391574 104614
rect 390954 68614 391574 104058
rect 390954 68058 390986 68614
rect 391542 68058 391574 68614
rect 390954 32614 391574 68058
rect 390954 32058 390986 32614
rect 391542 32058 391574 32614
rect 372954 -6662 372986 -6106
rect 373542 -6662 373574 -6106
rect 372954 -7654 373574 -6662
rect 390954 -7066 391574 32058
rect 397794 704838 398414 705830
rect 397794 704282 397826 704838
rect 398382 704282 398414 704838
rect 397794 687454 398414 704282
rect 397794 686898 397826 687454
rect 398382 686898 398414 687454
rect 397794 651454 398414 686898
rect 397794 650898 397826 651454
rect 398382 650898 398414 651454
rect 397794 615454 398414 650898
rect 397794 614898 397826 615454
rect 398382 614898 398414 615454
rect 397794 579454 398414 614898
rect 397794 578898 397826 579454
rect 398382 578898 398414 579454
rect 397794 543454 398414 578898
rect 397794 542898 397826 543454
rect 398382 542898 398414 543454
rect 397794 507454 398414 542898
rect 397794 506898 397826 507454
rect 398382 506898 398414 507454
rect 397794 471454 398414 506898
rect 397794 470898 397826 471454
rect 398382 470898 398414 471454
rect 397794 435454 398414 470898
rect 397794 434898 397826 435454
rect 398382 434898 398414 435454
rect 397794 399454 398414 434898
rect 397794 398898 397826 399454
rect 398382 398898 398414 399454
rect 397794 363454 398414 398898
rect 397794 362898 397826 363454
rect 398382 362898 398414 363454
rect 397794 327454 398414 362898
rect 397794 326898 397826 327454
rect 398382 326898 398414 327454
rect 397794 291454 398414 326898
rect 397794 290898 397826 291454
rect 398382 290898 398414 291454
rect 397794 255454 398414 290898
rect 397794 254898 397826 255454
rect 398382 254898 398414 255454
rect 397794 219454 398414 254898
rect 397794 218898 397826 219454
rect 398382 218898 398414 219454
rect 397794 183454 398414 218898
rect 397794 182898 397826 183454
rect 398382 182898 398414 183454
rect 397794 147454 398414 182898
rect 397794 146898 397826 147454
rect 398382 146898 398414 147454
rect 397794 111454 398414 146898
rect 397794 110898 397826 111454
rect 398382 110898 398414 111454
rect 397794 75454 398414 110898
rect 397794 74898 397826 75454
rect 398382 74898 398414 75454
rect 397794 39454 398414 74898
rect 397794 38898 397826 39454
rect 398382 38898 398414 39454
rect 397794 3454 398414 38898
rect 397794 2898 397826 3454
rect 398382 2898 398414 3454
rect 397794 -346 398414 2898
rect 397794 -902 397826 -346
rect 398382 -902 398414 -346
rect 397794 -1894 398414 -902
rect 401514 691174 402134 706202
rect 401514 690618 401546 691174
rect 402102 690618 402134 691174
rect 401514 655174 402134 690618
rect 401514 654618 401546 655174
rect 402102 654618 402134 655174
rect 401514 619174 402134 654618
rect 401514 618618 401546 619174
rect 402102 618618 402134 619174
rect 401514 583174 402134 618618
rect 401514 582618 401546 583174
rect 402102 582618 402134 583174
rect 401514 547174 402134 582618
rect 401514 546618 401546 547174
rect 402102 546618 402134 547174
rect 401514 511174 402134 546618
rect 401514 510618 401546 511174
rect 402102 510618 402134 511174
rect 401514 475174 402134 510618
rect 401514 474618 401546 475174
rect 402102 474618 402134 475174
rect 401514 439174 402134 474618
rect 401514 438618 401546 439174
rect 402102 438618 402134 439174
rect 401514 403174 402134 438618
rect 401514 402618 401546 403174
rect 402102 402618 402134 403174
rect 401514 367174 402134 402618
rect 401514 366618 401546 367174
rect 402102 366618 402134 367174
rect 401514 331174 402134 366618
rect 401514 330618 401546 331174
rect 402102 330618 402134 331174
rect 401514 295174 402134 330618
rect 401514 294618 401546 295174
rect 402102 294618 402134 295174
rect 401514 259174 402134 294618
rect 401514 258618 401546 259174
rect 402102 258618 402134 259174
rect 401514 223174 402134 258618
rect 401514 222618 401546 223174
rect 402102 222618 402134 223174
rect 401514 187174 402134 222618
rect 401514 186618 401546 187174
rect 402102 186618 402134 187174
rect 401514 151174 402134 186618
rect 401514 150618 401546 151174
rect 402102 150618 402134 151174
rect 401514 115174 402134 150618
rect 401514 114618 401546 115174
rect 402102 114618 402134 115174
rect 401514 79174 402134 114618
rect 401514 78618 401546 79174
rect 402102 78618 402134 79174
rect 401514 43174 402134 78618
rect 401514 42618 401546 43174
rect 402102 42618 402134 43174
rect 401514 7174 402134 42618
rect 401514 6618 401546 7174
rect 402102 6618 402134 7174
rect 401514 -2266 402134 6618
rect 401514 -2822 401546 -2266
rect 402102 -2822 402134 -2266
rect 401514 -3814 402134 -2822
rect 405234 694894 405854 708122
rect 405234 694338 405266 694894
rect 405822 694338 405854 694894
rect 405234 658894 405854 694338
rect 405234 658338 405266 658894
rect 405822 658338 405854 658894
rect 405234 622894 405854 658338
rect 405234 622338 405266 622894
rect 405822 622338 405854 622894
rect 405234 586894 405854 622338
rect 405234 586338 405266 586894
rect 405822 586338 405854 586894
rect 405234 550894 405854 586338
rect 405234 550338 405266 550894
rect 405822 550338 405854 550894
rect 405234 514894 405854 550338
rect 405234 514338 405266 514894
rect 405822 514338 405854 514894
rect 405234 478894 405854 514338
rect 405234 478338 405266 478894
rect 405822 478338 405854 478894
rect 405234 442894 405854 478338
rect 405234 442338 405266 442894
rect 405822 442338 405854 442894
rect 405234 406894 405854 442338
rect 405234 406338 405266 406894
rect 405822 406338 405854 406894
rect 405234 370894 405854 406338
rect 405234 370338 405266 370894
rect 405822 370338 405854 370894
rect 405234 334894 405854 370338
rect 405234 334338 405266 334894
rect 405822 334338 405854 334894
rect 405234 298894 405854 334338
rect 405234 298338 405266 298894
rect 405822 298338 405854 298894
rect 405234 262894 405854 298338
rect 405234 262338 405266 262894
rect 405822 262338 405854 262894
rect 405234 226894 405854 262338
rect 405234 226338 405266 226894
rect 405822 226338 405854 226894
rect 405234 190894 405854 226338
rect 405234 190338 405266 190894
rect 405822 190338 405854 190894
rect 405234 154894 405854 190338
rect 405234 154338 405266 154894
rect 405822 154338 405854 154894
rect 405234 118894 405854 154338
rect 405234 118338 405266 118894
rect 405822 118338 405854 118894
rect 405234 82894 405854 118338
rect 405234 82338 405266 82894
rect 405822 82338 405854 82894
rect 405234 46894 405854 82338
rect 405234 46338 405266 46894
rect 405822 46338 405854 46894
rect 405234 10894 405854 46338
rect 405234 10338 405266 10894
rect 405822 10338 405854 10894
rect 405234 -4186 405854 10338
rect 405234 -4742 405266 -4186
rect 405822 -4742 405854 -4186
rect 405234 -5734 405854 -4742
rect 408954 698614 409574 710042
rect 426954 711558 427574 711590
rect 426954 711002 426986 711558
rect 427542 711002 427574 711558
rect 423234 709638 423854 709670
rect 423234 709082 423266 709638
rect 423822 709082 423854 709638
rect 419514 707718 420134 707750
rect 419514 707162 419546 707718
rect 420102 707162 420134 707718
rect 408954 698058 408986 698614
rect 409542 698058 409574 698614
rect 408954 662614 409574 698058
rect 408954 662058 408986 662614
rect 409542 662058 409574 662614
rect 408954 626614 409574 662058
rect 408954 626058 408986 626614
rect 409542 626058 409574 626614
rect 408954 590614 409574 626058
rect 408954 590058 408986 590614
rect 409542 590058 409574 590614
rect 408954 554614 409574 590058
rect 408954 554058 408986 554614
rect 409542 554058 409574 554614
rect 408954 518614 409574 554058
rect 408954 518058 408986 518614
rect 409542 518058 409574 518614
rect 408954 482614 409574 518058
rect 408954 482058 408986 482614
rect 409542 482058 409574 482614
rect 408954 446614 409574 482058
rect 408954 446058 408986 446614
rect 409542 446058 409574 446614
rect 408954 410614 409574 446058
rect 408954 410058 408986 410614
rect 409542 410058 409574 410614
rect 408954 374614 409574 410058
rect 408954 374058 408986 374614
rect 409542 374058 409574 374614
rect 408954 338614 409574 374058
rect 408954 338058 408986 338614
rect 409542 338058 409574 338614
rect 408954 302614 409574 338058
rect 408954 302058 408986 302614
rect 409542 302058 409574 302614
rect 408954 266614 409574 302058
rect 408954 266058 408986 266614
rect 409542 266058 409574 266614
rect 408954 230614 409574 266058
rect 408954 230058 408986 230614
rect 409542 230058 409574 230614
rect 408954 194614 409574 230058
rect 408954 194058 408986 194614
rect 409542 194058 409574 194614
rect 408954 158614 409574 194058
rect 408954 158058 408986 158614
rect 409542 158058 409574 158614
rect 408954 122614 409574 158058
rect 408954 122058 408986 122614
rect 409542 122058 409574 122614
rect 408954 86614 409574 122058
rect 408954 86058 408986 86614
rect 409542 86058 409574 86614
rect 408954 50614 409574 86058
rect 408954 50058 408986 50614
rect 409542 50058 409574 50614
rect 408954 14614 409574 50058
rect 408954 14058 408986 14614
rect 409542 14058 409574 14614
rect 390954 -7622 390986 -7066
rect 391542 -7622 391574 -7066
rect 390954 -7654 391574 -7622
rect 408954 -6106 409574 14058
rect 415794 705798 416414 705830
rect 415794 705242 415826 705798
rect 416382 705242 416414 705798
rect 415794 669454 416414 705242
rect 415794 668898 415826 669454
rect 416382 668898 416414 669454
rect 415794 633454 416414 668898
rect 415794 632898 415826 633454
rect 416382 632898 416414 633454
rect 415794 597454 416414 632898
rect 415794 596898 415826 597454
rect 416382 596898 416414 597454
rect 415794 561454 416414 596898
rect 415794 560898 415826 561454
rect 416382 560898 416414 561454
rect 415794 525454 416414 560898
rect 415794 524898 415826 525454
rect 416382 524898 416414 525454
rect 415794 489454 416414 524898
rect 415794 488898 415826 489454
rect 416382 488898 416414 489454
rect 415794 453454 416414 488898
rect 415794 452898 415826 453454
rect 416382 452898 416414 453454
rect 415794 417454 416414 452898
rect 415794 416898 415826 417454
rect 416382 416898 416414 417454
rect 415794 381454 416414 416898
rect 415794 380898 415826 381454
rect 416382 380898 416414 381454
rect 415794 345454 416414 380898
rect 415794 344898 415826 345454
rect 416382 344898 416414 345454
rect 415794 309454 416414 344898
rect 415794 308898 415826 309454
rect 416382 308898 416414 309454
rect 415794 273454 416414 308898
rect 415794 272898 415826 273454
rect 416382 272898 416414 273454
rect 415794 237454 416414 272898
rect 415794 236898 415826 237454
rect 416382 236898 416414 237454
rect 415794 201454 416414 236898
rect 415794 200898 415826 201454
rect 416382 200898 416414 201454
rect 415794 165454 416414 200898
rect 415794 164898 415826 165454
rect 416382 164898 416414 165454
rect 415794 129454 416414 164898
rect 415794 128898 415826 129454
rect 416382 128898 416414 129454
rect 415794 93454 416414 128898
rect 415794 92898 415826 93454
rect 416382 92898 416414 93454
rect 415794 57454 416414 92898
rect 415794 56898 415826 57454
rect 416382 56898 416414 57454
rect 415794 21454 416414 56898
rect 415794 20898 415826 21454
rect 416382 20898 416414 21454
rect 415794 -1306 416414 20898
rect 415794 -1862 415826 -1306
rect 416382 -1862 416414 -1306
rect 415794 -1894 416414 -1862
rect 419514 673174 420134 707162
rect 419514 672618 419546 673174
rect 420102 672618 420134 673174
rect 419514 637174 420134 672618
rect 419514 636618 419546 637174
rect 420102 636618 420134 637174
rect 419514 601174 420134 636618
rect 419514 600618 419546 601174
rect 420102 600618 420134 601174
rect 419514 565174 420134 600618
rect 419514 564618 419546 565174
rect 420102 564618 420134 565174
rect 419514 529174 420134 564618
rect 419514 528618 419546 529174
rect 420102 528618 420134 529174
rect 419514 493174 420134 528618
rect 419514 492618 419546 493174
rect 420102 492618 420134 493174
rect 419514 457174 420134 492618
rect 419514 456618 419546 457174
rect 420102 456618 420134 457174
rect 419514 421174 420134 456618
rect 419514 420618 419546 421174
rect 420102 420618 420134 421174
rect 419514 385174 420134 420618
rect 419514 384618 419546 385174
rect 420102 384618 420134 385174
rect 419514 349174 420134 384618
rect 419514 348618 419546 349174
rect 420102 348618 420134 349174
rect 419514 313174 420134 348618
rect 419514 312618 419546 313174
rect 420102 312618 420134 313174
rect 419514 277174 420134 312618
rect 419514 276618 419546 277174
rect 420102 276618 420134 277174
rect 419514 241174 420134 276618
rect 419514 240618 419546 241174
rect 420102 240618 420134 241174
rect 419514 205174 420134 240618
rect 419514 204618 419546 205174
rect 420102 204618 420134 205174
rect 419514 169174 420134 204618
rect 419514 168618 419546 169174
rect 420102 168618 420134 169174
rect 419514 133174 420134 168618
rect 419514 132618 419546 133174
rect 420102 132618 420134 133174
rect 419514 97174 420134 132618
rect 419514 96618 419546 97174
rect 420102 96618 420134 97174
rect 419514 61174 420134 96618
rect 419514 60618 419546 61174
rect 420102 60618 420134 61174
rect 419514 25174 420134 60618
rect 419514 24618 419546 25174
rect 420102 24618 420134 25174
rect 419514 -3226 420134 24618
rect 419514 -3782 419546 -3226
rect 420102 -3782 420134 -3226
rect 419514 -3814 420134 -3782
rect 423234 676894 423854 709082
rect 423234 676338 423266 676894
rect 423822 676338 423854 676894
rect 423234 640894 423854 676338
rect 423234 640338 423266 640894
rect 423822 640338 423854 640894
rect 423234 604894 423854 640338
rect 423234 604338 423266 604894
rect 423822 604338 423854 604894
rect 423234 568894 423854 604338
rect 423234 568338 423266 568894
rect 423822 568338 423854 568894
rect 423234 532894 423854 568338
rect 423234 532338 423266 532894
rect 423822 532338 423854 532894
rect 423234 496894 423854 532338
rect 423234 496338 423266 496894
rect 423822 496338 423854 496894
rect 423234 460894 423854 496338
rect 423234 460338 423266 460894
rect 423822 460338 423854 460894
rect 423234 424894 423854 460338
rect 423234 424338 423266 424894
rect 423822 424338 423854 424894
rect 423234 388894 423854 424338
rect 423234 388338 423266 388894
rect 423822 388338 423854 388894
rect 423234 352894 423854 388338
rect 423234 352338 423266 352894
rect 423822 352338 423854 352894
rect 423234 316894 423854 352338
rect 423234 316338 423266 316894
rect 423822 316338 423854 316894
rect 423234 280894 423854 316338
rect 423234 280338 423266 280894
rect 423822 280338 423854 280894
rect 423234 244894 423854 280338
rect 423234 244338 423266 244894
rect 423822 244338 423854 244894
rect 423234 208894 423854 244338
rect 423234 208338 423266 208894
rect 423822 208338 423854 208894
rect 423234 172894 423854 208338
rect 423234 172338 423266 172894
rect 423822 172338 423854 172894
rect 423234 136894 423854 172338
rect 423234 136338 423266 136894
rect 423822 136338 423854 136894
rect 423234 100894 423854 136338
rect 423234 100338 423266 100894
rect 423822 100338 423854 100894
rect 423234 64894 423854 100338
rect 423234 64338 423266 64894
rect 423822 64338 423854 64894
rect 423234 28894 423854 64338
rect 423234 28338 423266 28894
rect 423822 28338 423854 28894
rect 423234 -5146 423854 28338
rect 423234 -5702 423266 -5146
rect 423822 -5702 423854 -5146
rect 423234 -5734 423854 -5702
rect 426954 680614 427574 711002
rect 444954 710598 445574 711590
rect 444954 710042 444986 710598
rect 445542 710042 445574 710598
rect 441234 708678 441854 709670
rect 441234 708122 441266 708678
rect 441822 708122 441854 708678
rect 437514 706758 438134 707750
rect 437514 706202 437546 706758
rect 438102 706202 438134 706758
rect 426954 680058 426986 680614
rect 427542 680058 427574 680614
rect 426954 644614 427574 680058
rect 426954 644058 426986 644614
rect 427542 644058 427574 644614
rect 426954 608614 427574 644058
rect 426954 608058 426986 608614
rect 427542 608058 427574 608614
rect 426954 572614 427574 608058
rect 426954 572058 426986 572614
rect 427542 572058 427574 572614
rect 426954 536614 427574 572058
rect 426954 536058 426986 536614
rect 427542 536058 427574 536614
rect 426954 500614 427574 536058
rect 426954 500058 426986 500614
rect 427542 500058 427574 500614
rect 426954 464614 427574 500058
rect 426954 464058 426986 464614
rect 427542 464058 427574 464614
rect 426954 428614 427574 464058
rect 426954 428058 426986 428614
rect 427542 428058 427574 428614
rect 426954 392614 427574 428058
rect 426954 392058 426986 392614
rect 427542 392058 427574 392614
rect 426954 356614 427574 392058
rect 426954 356058 426986 356614
rect 427542 356058 427574 356614
rect 426954 320614 427574 356058
rect 426954 320058 426986 320614
rect 427542 320058 427574 320614
rect 426954 284614 427574 320058
rect 426954 284058 426986 284614
rect 427542 284058 427574 284614
rect 426954 248614 427574 284058
rect 426954 248058 426986 248614
rect 427542 248058 427574 248614
rect 426954 212614 427574 248058
rect 426954 212058 426986 212614
rect 427542 212058 427574 212614
rect 426954 176614 427574 212058
rect 426954 176058 426986 176614
rect 427542 176058 427574 176614
rect 426954 140614 427574 176058
rect 426954 140058 426986 140614
rect 427542 140058 427574 140614
rect 426954 104614 427574 140058
rect 426954 104058 426986 104614
rect 427542 104058 427574 104614
rect 426954 68614 427574 104058
rect 426954 68058 426986 68614
rect 427542 68058 427574 68614
rect 426954 32614 427574 68058
rect 426954 32058 426986 32614
rect 427542 32058 427574 32614
rect 408954 -6662 408986 -6106
rect 409542 -6662 409574 -6106
rect 408954 -7654 409574 -6662
rect 426954 -7066 427574 32058
rect 433794 704838 434414 705830
rect 433794 704282 433826 704838
rect 434382 704282 434414 704838
rect 433794 687454 434414 704282
rect 433794 686898 433826 687454
rect 434382 686898 434414 687454
rect 433794 651454 434414 686898
rect 433794 650898 433826 651454
rect 434382 650898 434414 651454
rect 433794 615454 434414 650898
rect 433794 614898 433826 615454
rect 434382 614898 434414 615454
rect 433794 579454 434414 614898
rect 433794 578898 433826 579454
rect 434382 578898 434414 579454
rect 433794 543454 434414 578898
rect 433794 542898 433826 543454
rect 434382 542898 434414 543454
rect 433794 507454 434414 542898
rect 433794 506898 433826 507454
rect 434382 506898 434414 507454
rect 433794 471454 434414 506898
rect 433794 470898 433826 471454
rect 434382 470898 434414 471454
rect 433794 435454 434414 470898
rect 433794 434898 433826 435454
rect 434382 434898 434414 435454
rect 433794 399454 434414 434898
rect 433794 398898 433826 399454
rect 434382 398898 434414 399454
rect 433794 363454 434414 398898
rect 433794 362898 433826 363454
rect 434382 362898 434414 363454
rect 433794 327454 434414 362898
rect 433794 326898 433826 327454
rect 434382 326898 434414 327454
rect 433794 291454 434414 326898
rect 433794 290898 433826 291454
rect 434382 290898 434414 291454
rect 433794 255454 434414 290898
rect 433794 254898 433826 255454
rect 434382 254898 434414 255454
rect 433794 219454 434414 254898
rect 433794 218898 433826 219454
rect 434382 218898 434414 219454
rect 433794 183454 434414 218898
rect 433794 182898 433826 183454
rect 434382 182898 434414 183454
rect 433794 147454 434414 182898
rect 433794 146898 433826 147454
rect 434382 146898 434414 147454
rect 433794 111454 434414 146898
rect 433794 110898 433826 111454
rect 434382 110898 434414 111454
rect 433794 75454 434414 110898
rect 433794 74898 433826 75454
rect 434382 74898 434414 75454
rect 433794 39454 434414 74898
rect 433794 38898 433826 39454
rect 434382 38898 434414 39454
rect 433794 3454 434414 38898
rect 433794 2898 433826 3454
rect 434382 2898 434414 3454
rect 433794 -346 434414 2898
rect 433794 -902 433826 -346
rect 434382 -902 434414 -346
rect 433794 -1894 434414 -902
rect 437514 691174 438134 706202
rect 437514 690618 437546 691174
rect 438102 690618 438134 691174
rect 437514 655174 438134 690618
rect 437514 654618 437546 655174
rect 438102 654618 438134 655174
rect 437514 619174 438134 654618
rect 437514 618618 437546 619174
rect 438102 618618 438134 619174
rect 437514 583174 438134 618618
rect 437514 582618 437546 583174
rect 438102 582618 438134 583174
rect 437514 547174 438134 582618
rect 437514 546618 437546 547174
rect 438102 546618 438134 547174
rect 437514 511174 438134 546618
rect 437514 510618 437546 511174
rect 438102 510618 438134 511174
rect 437514 475174 438134 510618
rect 437514 474618 437546 475174
rect 438102 474618 438134 475174
rect 437514 439174 438134 474618
rect 437514 438618 437546 439174
rect 438102 438618 438134 439174
rect 437514 403174 438134 438618
rect 437514 402618 437546 403174
rect 438102 402618 438134 403174
rect 437514 367174 438134 402618
rect 437514 366618 437546 367174
rect 438102 366618 438134 367174
rect 437514 331174 438134 366618
rect 437514 330618 437546 331174
rect 438102 330618 438134 331174
rect 437514 295174 438134 330618
rect 437514 294618 437546 295174
rect 438102 294618 438134 295174
rect 437514 259174 438134 294618
rect 437514 258618 437546 259174
rect 438102 258618 438134 259174
rect 437514 223174 438134 258618
rect 437514 222618 437546 223174
rect 438102 222618 438134 223174
rect 437514 187174 438134 222618
rect 437514 186618 437546 187174
rect 438102 186618 438134 187174
rect 437514 151174 438134 186618
rect 437514 150618 437546 151174
rect 438102 150618 438134 151174
rect 437514 115174 438134 150618
rect 437514 114618 437546 115174
rect 438102 114618 438134 115174
rect 437514 79174 438134 114618
rect 437514 78618 437546 79174
rect 438102 78618 438134 79174
rect 437514 43174 438134 78618
rect 437514 42618 437546 43174
rect 438102 42618 438134 43174
rect 437514 7174 438134 42618
rect 437514 6618 437546 7174
rect 438102 6618 438134 7174
rect 437514 -2266 438134 6618
rect 437514 -2822 437546 -2266
rect 438102 -2822 438134 -2266
rect 437514 -3814 438134 -2822
rect 441234 694894 441854 708122
rect 441234 694338 441266 694894
rect 441822 694338 441854 694894
rect 441234 658894 441854 694338
rect 441234 658338 441266 658894
rect 441822 658338 441854 658894
rect 441234 622894 441854 658338
rect 441234 622338 441266 622894
rect 441822 622338 441854 622894
rect 441234 586894 441854 622338
rect 441234 586338 441266 586894
rect 441822 586338 441854 586894
rect 441234 550894 441854 586338
rect 441234 550338 441266 550894
rect 441822 550338 441854 550894
rect 441234 514894 441854 550338
rect 441234 514338 441266 514894
rect 441822 514338 441854 514894
rect 441234 478894 441854 514338
rect 441234 478338 441266 478894
rect 441822 478338 441854 478894
rect 441234 442894 441854 478338
rect 441234 442338 441266 442894
rect 441822 442338 441854 442894
rect 441234 406894 441854 442338
rect 441234 406338 441266 406894
rect 441822 406338 441854 406894
rect 441234 370894 441854 406338
rect 441234 370338 441266 370894
rect 441822 370338 441854 370894
rect 441234 334894 441854 370338
rect 441234 334338 441266 334894
rect 441822 334338 441854 334894
rect 441234 298894 441854 334338
rect 441234 298338 441266 298894
rect 441822 298338 441854 298894
rect 441234 262894 441854 298338
rect 441234 262338 441266 262894
rect 441822 262338 441854 262894
rect 441234 226894 441854 262338
rect 441234 226338 441266 226894
rect 441822 226338 441854 226894
rect 441234 190894 441854 226338
rect 441234 190338 441266 190894
rect 441822 190338 441854 190894
rect 441234 154894 441854 190338
rect 441234 154338 441266 154894
rect 441822 154338 441854 154894
rect 441234 118894 441854 154338
rect 441234 118338 441266 118894
rect 441822 118338 441854 118894
rect 441234 82894 441854 118338
rect 441234 82338 441266 82894
rect 441822 82338 441854 82894
rect 441234 46894 441854 82338
rect 441234 46338 441266 46894
rect 441822 46338 441854 46894
rect 441234 10894 441854 46338
rect 441234 10338 441266 10894
rect 441822 10338 441854 10894
rect 441234 -4186 441854 10338
rect 441234 -4742 441266 -4186
rect 441822 -4742 441854 -4186
rect 441234 -5734 441854 -4742
rect 444954 698614 445574 710042
rect 462954 711558 463574 711590
rect 462954 711002 462986 711558
rect 463542 711002 463574 711558
rect 459234 709638 459854 709670
rect 459234 709082 459266 709638
rect 459822 709082 459854 709638
rect 455514 707718 456134 707750
rect 455514 707162 455546 707718
rect 456102 707162 456134 707718
rect 444954 698058 444986 698614
rect 445542 698058 445574 698614
rect 444954 662614 445574 698058
rect 444954 662058 444986 662614
rect 445542 662058 445574 662614
rect 444954 626614 445574 662058
rect 444954 626058 444986 626614
rect 445542 626058 445574 626614
rect 444954 590614 445574 626058
rect 444954 590058 444986 590614
rect 445542 590058 445574 590614
rect 444954 554614 445574 590058
rect 444954 554058 444986 554614
rect 445542 554058 445574 554614
rect 444954 518614 445574 554058
rect 444954 518058 444986 518614
rect 445542 518058 445574 518614
rect 444954 482614 445574 518058
rect 444954 482058 444986 482614
rect 445542 482058 445574 482614
rect 444954 446614 445574 482058
rect 444954 446058 444986 446614
rect 445542 446058 445574 446614
rect 444954 410614 445574 446058
rect 444954 410058 444986 410614
rect 445542 410058 445574 410614
rect 444954 374614 445574 410058
rect 444954 374058 444986 374614
rect 445542 374058 445574 374614
rect 444954 338614 445574 374058
rect 444954 338058 444986 338614
rect 445542 338058 445574 338614
rect 444954 302614 445574 338058
rect 444954 302058 444986 302614
rect 445542 302058 445574 302614
rect 444954 266614 445574 302058
rect 444954 266058 444986 266614
rect 445542 266058 445574 266614
rect 444954 230614 445574 266058
rect 444954 230058 444986 230614
rect 445542 230058 445574 230614
rect 444954 194614 445574 230058
rect 444954 194058 444986 194614
rect 445542 194058 445574 194614
rect 444954 158614 445574 194058
rect 444954 158058 444986 158614
rect 445542 158058 445574 158614
rect 444954 122614 445574 158058
rect 444954 122058 444986 122614
rect 445542 122058 445574 122614
rect 444954 86614 445574 122058
rect 444954 86058 444986 86614
rect 445542 86058 445574 86614
rect 444954 50614 445574 86058
rect 444954 50058 444986 50614
rect 445542 50058 445574 50614
rect 444954 14614 445574 50058
rect 444954 14058 444986 14614
rect 445542 14058 445574 14614
rect 426954 -7622 426986 -7066
rect 427542 -7622 427574 -7066
rect 426954 -7654 427574 -7622
rect 444954 -6106 445574 14058
rect 451794 705798 452414 705830
rect 451794 705242 451826 705798
rect 452382 705242 452414 705798
rect 451794 669454 452414 705242
rect 451794 668898 451826 669454
rect 452382 668898 452414 669454
rect 451794 633454 452414 668898
rect 451794 632898 451826 633454
rect 452382 632898 452414 633454
rect 451794 597454 452414 632898
rect 451794 596898 451826 597454
rect 452382 596898 452414 597454
rect 451794 561454 452414 596898
rect 451794 560898 451826 561454
rect 452382 560898 452414 561454
rect 451794 525454 452414 560898
rect 451794 524898 451826 525454
rect 452382 524898 452414 525454
rect 451794 489454 452414 524898
rect 451794 488898 451826 489454
rect 452382 488898 452414 489454
rect 451794 453454 452414 488898
rect 451794 452898 451826 453454
rect 452382 452898 452414 453454
rect 451794 417454 452414 452898
rect 451794 416898 451826 417454
rect 452382 416898 452414 417454
rect 451794 381454 452414 416898
rect 451794 380898 451826 381454
rect 452382 380898 452414 381454
rect 451794 345454 452414 380898
rect 451794 344898 451826 345454
rect 452382 344898 452414 345454
rect 451794 309454 452414 344898
rect 451794 308898 451826 309454
rect 452382 308898 452414 309454
rect 451794 273454 452414 308898
rect 451794 272898 451826 273454
rect 452382 272898 452414 273454
rect 451794 237454 452414 272898
rect 451794 236898 451826 237454
rect 452382 236898 452414 237454
rect 451794 201454 452414 236898
rect 451794 200898 451826 201454
rect 452382 200898 452414 201454
rect 451794 165454 452414 200898
rect 451794 164898 451826 165454
rect 452382 164898 452414 165454
rect 451794 129454 452414 164898
rect 451794 128898 451826 129454
rect 452382 128898 452414 129454
rect 451794 93454 452414 128898
rect 451794 92898 451826 93454
rect 452382 92898 452414 93454
rect 451794 57454 452414 92898
rect 451794 56898 451826 57454
rect 452382 56898 452414 57454
rect 451794 21454 452414 56898
rect 451794 20898 451826 21454
rect 452382 20898 452414 21454
rect 451794 -1306 452414 20898
rect 451794 -1862 451826 -1306
rect 452382 -1862 452414 -1306
rect 451794 -1894 452414 -1862
rect 455514 673174 456134 707162
rect 455514 672618 455546 673174
rect 456102 672618 456134 673174
rect 455514 637174 456134 672618
rect 455514 636618 455546 637174
rect 456102 636618 456134 637174
rect 455514 601174 456134 636618
rect 455514 600618 455546 601174
rect 456102 600618 456134 601174
rect 455514 565174 456134 600618
rect 455514 564618 455546 565174
rect 456102 564618 456134 565174
rect 455514 529174 456134 564618
rect 455514 528618 455546 529174
rect 456102 528618 456134 529174
rect 455514 493174 456134 528618
rect 455514 492618 455546 493174
rect 456102 492618 456134 493174
rect 455514 457174 456134 492618
rect 455514 456618 455546 457174
rect 456102 456618 456134 457174
rect 455514 421174 456134 456618
rect 455514 420618 455546 421174
rect 456102 420618 456134 421174
rect 455514 385174 456134 420618
rect 455514 384618 455546 385174
rect 456102 384618 456134 385174
rect 455514 349174 456134 384618
rect 455514 348618 455546 349174
rect 456102 348618 456134 349174
rect 455514 313174 456134 348618
rect 455514 312618 455546 313174
rect 456102 312618 456134 313174
rect 455514 277174 456134 312618
rect 455514 276618 455546 277174
rect 456102 276618 456134 277174
rect 455514 241174 456134 276618
rect 455514 240618 455546 241174
rect 456102 240618 456134 241174
rect 455514 205174 456134 240618
rect 455514 204618 455546 205174
rect 456102 204618 456134 205174
rect 455514 169174 456134 204618
rect 455514 168618 455546 169174
rect 456102 168618 456134 169174
rect 455514 133174 456134 168618
rect 455514 132618 455546 133174
rect 456102 132618 456134 133174
rect 455514 97174 456134 132618
rect 455514 96618 455546 97174
rect 456102 96618 456134 97174
rect 455514 61174 456134 96618
rect 455514 60618 455546 61174
rect 456102 60618 456134 61174
rect 455514 25174 456134 60618
rect 455514 24618 455546 25174
rect 456102 24618 456134 25174
rect 455514 -3226 456134 24618
rect 455514 -3782 455546 -3226
rect 456102 -3782 456134 -3226
rect 455514 -3814 456134 -3782
rect 459234 676894 459854 709082
rect 459234 676338 459266 676894
rect 459822 676338 459854 676894
rect 459234 640894 459854 676338
rect 459234 640338 459266 640894
rect 459822 640338 459854 640894
rect 459234 604894 459854 640338
rect 459234 604338 459266 604894
rect 459822 604338 459854 604894
rect 459234 568894 459854 604338
rect 459234 568338 459266 568894
rect 459822 568338 459854 568894
rect 459234 532894 459854 568338
rect 459234 532338 459266 532894
rect 459822 532338 459854 532894
rect 459234 496894 459854 532338
rect 459234 496338 459266 496894
rect 459822 496338 459854 496894
rect 459234 460894 459854 496338
rect 459234 460338 459266 460894
rect 459822 460338 459854 460894
rect 459234 424894 459854 460338
rect 459234 424338 459266 424894
rect 459822 424338 459854 424894
rect 459234 388894 459854 424338
rect 459234 388338 459266 388894
rect 459822 388338 459854 388894
rect 459234 352894 459854 388338
rect 459234 352338 459266 352894
rect 459822 352338 459854 352894
rect 459234 316894 459854 352338
rect 459234 316338 459266 316894
rect 459822 316338 459854 316894
rect 459234 280894 459854 316338
rect 459234 280338 459266 280894
rect 459822 280338 459854 280894
rect 459234 244894 459854 280338
rect 459234 244338 459266 244894
rect 459822 244338 459854 244894
rect 459234 208894 459854 244338
rect 459234 208338 459266 208894
rect 459822 208338 459854 208894
rect 459234 172894 459854 208338
rect 459234 172338 459266 172894
rect 459822 172338 459854 172894
rect 459234 136894 459854 172338
rect 459234 136338 459266 136894
rect 459822 136338 459854 136894
rect 459234 100894 459854 136338
rect 459234 100338 459266 100894
rect 459822 100338 459854 100894
rect 459234 64894 459854 100338
rect 459234 64338 459266 64894
rect 459822 64338 459854 64894
rect 459234 28894 459854 64338
rect 459234 28338 459266 28894
rect 459822 28338 459854 28894
rect 459234 -5146 459854 28338
rect 459234 -5702 459266 -5146
rect 459822 -5702 459854 -5146
rect 459234 -5734 459854 -5702
rect 462954 680614 463574 711002
rect 480954 710598 481574 711590
rect 480954 710042 480986 710598
rect 481542 710042 481574 710598
rect 477234 708678 477854 709670
rect 477234 708122 477266 708678
rect 477822 708122 477854 708678
rect 473514 706758 474134 707750
rect 473514 706202 473546 706758
rect 474102 706202 474134 706758
rect 462954 680058 462986 680614
rect 463542 680058 463574 680614
rect 462954 644614 463574 680058
rect 462954 644058 462986 644614
rect 463542 644058 463574 644614
rect 462954 608614 463574 644058
rect 462954 608058 462986 608614
rect 463542 608058 463574 608614
rect 462954 572614 463574 608058
rect 462954 572058 462986 572614
rect 463542 572058 463574 572614
rect 462954 536614 463574 572058
rect 462954 536058 462986 536614
rect 463542 536058 463574 536614
rect 462954 500614 463574 536058
rect 462954 500058 462986 500614
rect 463542 500058 463574 500614
rect 462954 464614 463574 500058
rect 462954 464058 462986 464614
rect 463542 464058 463574 464614
rect 462954 428614 463574 464058
rect 462954 428058 462986 428614
rect 463542 428058 463574 428614
rect 462954 392614 463574 428058
rect 462954 392058 462986 392614
rect 463542 392058 463574 392614
rect 462954 356614 463574 392058
rect 462954 356058 462986 356614
rect 463542 356058 463574 356614
rect 462954 320614 463574 356058
rect 462954 320058 462986 320614
rect 463542 320058 463574 320614
rect 462954 284614 463574 320058
rect 462954 284058 462986 284614
rect 463542 284058 463574 284614
rect 462954 248614 463574 284058
rect 462954 248058 462986 248614
rect 463542 248058 463574 248614
rect 462954 212614 463574 248058
rect 462954 212058 462986 212614
rect 463542 212058 463574 212614
rect 462954 176614 463574 212058
rect 462954 176058 462986 176614
rect 463542 176058 463574 176614
rect 462954 140614 463574 176058
rect 462954 140058 462986 140614
rect 463542 140058 463574 140614
rect 462954 104614 463574 140058
rect 462954 104058 462986 104614
rect 463542 104058 463574 104614
rect 462954 68614 463574 104058
rect 462954 68058 462986 68614
rect 463542 68058 463574 68614
rect 462954 32614 463574 68058
rect 462954 32058 462986 32614
rect 463542 32058 463574 32614
rect 444954 -6662 444986 -6106
rect 445542 -6662 445574 -6106
rect 444954 -7654 445574 -6662
rect 462954 -7066 463574 32058
rect 469794 704838 470414 705830
rect 469794 704282 469826 704838
rect 470382 704282 470414 704838
rect 469794 687454 470414 704282
rect 469794 686898 469826 687454
rect 470382 686898 470414 687454
rect 469794 651454 470414 686898
rect 469794 650898 469826 651454
rect 470382 650898 470414 651454
rect 469794 615454 470414 650898
rect 469794 614898 469826 615454
rect 470382 614898 470414 615454
rect 469794 579454 470414 614898
rect 469794 578898 469826 579454
rect 470382 578898 470414 579454
rect 469794 543454 470414 578898
rect 469794 542898 469826 543454
rect 470382 542898 470414 543454
rect 469794 507454 470414 542898
rect 469794 506898 469826 507454
rect 470382 506898 470414 507454
rect 469794 471454 470414 506898
rect 469794 470898 469826 471454
rect 470382 470898 470414 471454
rect 469794 435454 470414 470898
rect 469794 434898 469826 435454
rect 470382 434898 470414 435454
rect 469794 399454 470414 434898
rect 469794 398898 469826 399454
rect 470382 398898 470414 399454
rect 469794 363454 470414 398898
rect 469794 362898 469826 363454
rect 470382 362898 470414 363454
rect 469794 327454 470414 362898
rect 469794 326898 469826 327454
rect 470382 326898 470414 327454
rect 469794 291454 470414 326898
rect 469794 290898 469826 291454
rect 470382 290898 470414 291454
rect 469794 255454 470414 290898
rect 469794 254898 469826 255454
rect 470382 254898 470414 255454
rect 469794 219454 470414 254898
rect 469794 218898 469826 219454
rect 470382 218898 470414 219454
rect 469794 183454 470414 218898
rect 469794 182898 469826 183454
rect 470382 182898 470414 183454
rect 469794 147454 470414 182898
rect 469794 146898 469826 147454
rect 470382 146898 470414 147454
rect 469794 111454 470414 146898
rect 469794 110898 469826 111454
rect 470382 110898 470414 111454
rect 469794 75454 470414 110898
rect 469794 74898 469826 75454
rect 470382 74898 470414 75454
rect 469794 39454 470414 74898
rect 469794 38898 469826 39454
rect 470382 38898 470414 39454
rect 469794 3454 470414 38898
rect 469794 2898 469826 3454
rect 470382 2898 470414 3454
rect 469794 -346 470414 2898
rect 469794 -902 469826 -346
rect 470382 -902 470414 -346
rect 469794 -1894 470414 -902
rect 473514 691174 474134 706202
rect 473514 690618 473546 691174
rect 474102 690618 474134 691174
rect 473514 655174 474134 690618
rect 473514 654618 473546 655174
rect 474102 654618 474134 655174
rect 473514 619174 474134 654618
rect 473514 618618 473546 619174
rect 474102 618618 474134 619174
rect 473514 583174 474134 618618
rect 473514 582618 473546 583174
rect 474102 582618 474134 583174
rect 473514 547174 474134 582618
rect 473514 546618 473546 547174
rect 474102 546618 474134 547174
rect 473514 511174 474134 546618
rect 473514 510618 473546 511174
rect 474102 510618 474134 511174
rect 473514 475174 474134 510618
rect 473514 474618 473546 475174
rect 474102 474618 474134 475174
rect 473514 439174 474134 474618
rect 473514 438618 473546 439174
rect 474102 438618 474134 439174
rect 473514 403174 474134 438618
rect 473514 402618 473546 403174
rect 474102 402618 474134 403174
rect 473514 367174 474134 402618
rect 473514 366618 473546 367174
rect 474102 366618 474134 367174
rect 473514 331174 474134 366618
rect 473514 330618 473546 331174
rect 474102 330618 474134 331174
rect 473514 295174 474134 330618
rect 473514 294618 473546 295174
rect 474102 294618 474134 295174
rect 473514 259174 474134 294618
rect 473514 258618 473546 259174
rect 474102 258618 474134 259174
rect 473514 223174 474134 258618
rect 473514 222618 473546 223174
rect 474102 222618 474134 223174
rect 473514 187174 474134 222618
rect 473514 186618 473546 187174
rect 474102 186618 474134 187174
rect 473514 151174 474134 186618
rect 473514 150618 473546 151174
rect 474102 150618 474134 151174
rect 473514 115174 474134 150618
rect 473514 114618 473546 115174
rect 474102 114618 474134 115174
rect 473514 79174 474134 114618
rect 473514 78618 473546 79174
rect 474102 78618 474134 79174
rect 473514 43174 474134 78618
rect 473514 42618 473546 43174
rect 474102 42618 474134 43174
rect 473514 7174 474134 42618
rect 473514 6618 473546 7174
rect 474102 6618 474134 7174
rect 473514 -2266 474134 6618
rect 473514 -2822 473546 -2266
rect 474102 -2822 474134 -2266
rect 473514 -3814 474134 -2822
rect 477234 694894 477854 708122
rect 477234 694338 477266 694894
rect 477822 694338 477854 694894
rect 477234 658894 477854 694338
rect 477234 658338 477266 658894
rect 477822 658338 477854 658894
rect 477234 622894 477854 658338
rect 477234 622338 477266 622894
rect 477822 622338 477854 622894
rect 477234 586894 477854 622338
rect 477234 586338 477266 586894
rect 477822 586338 477854 586894
rect 477234 550894 477854 586338
rect 477234 550338 477266 550894
rect 477822 550338 477854 550894
rect 477234 514894 477854 550338
rect 477234 514338 477266 514894
rect 477822 514338 477854 514894
rect 477234 478894 477854 514338
rect 477234 478338 477266 478894
rect 477822 478338 477854 478894
rect 477234 442894 477854 478338
rect 477234 442338 477266 442894
rect 477822 442338 477854 442894
rect 477234 406894 477854 442338
rect 477234 406338 477266 406894
rect 477822 406338 477854 406894
rect 477234 370894 477854 406338
rect 477234 370338 477266 370894
rect 477822 370338 477854 370894
rect 477234 334894 477854 370338
rect 477234 334338 477266 334894
rect 477822 334338 477854 334894
rect 477234 298894 477854 334338
rect 477234 298338 477266 298894
rect 477822 298338 477854 298894
rect 477234 262894 477854 298338
rect 477234 262338 477266 262894
rect 477822 262338 477854 262894
rect 477234 226894 477854 262338
rect 477234 226338 477266 226894
rect 477822 226338 477854 226894
rect 477234 190894 477854 226338
rect 477234 190338 477266 190894
rect 477822 190338 477854 190894
rect 477234 154894 477854 190338
rect 477234 154338 477266 154894
rect 477822 154338 477854 154894
rect 477234 118894 477854 154338
rect 477234 118338 477266 118894
rect 477822 118338 477854 118894
rect 477234 82894 477854 118338
rect 477234 82338 477266 82894
rect 477822 82338 477854 82894
rect 477234 46894 477854 82338
rect 477234 46338 477266 46894
rect 477822 46338 477854 46894
rect 477234 10894 477854 46338
rect 477234 10338 477266 10894
rect 477822 10338 477854 10894
rect 477234 -4186 477854 10338
rect 477234 -4742 477266 -4186
rect 477822 -4742 477854 -4186
rect 477234 -5734 477854 -4742
rect 480954 698614 481574 710042
rect 498954 711558 499574 711590
rect 498954 711002 498986 711558
rect 499542 711002 499574 711558
rect 495234 709638 495854 709670
rect 495234 709082 495266 709638
rect 495822 709082 495854 709638
rect 491514 707718 492134 707750
rect 491514 707162 491546 707718
rect 492102 707162 492134 707718
rect 480954 698058 480986 698614
rect 481542 698058 481574 698614
rect 480954 662614 481574 698058
rect 480954 662058 480986 662614
rect 481542 662058 481574 662614
rect 480954 626614 481574 662058
rect 480954 626058 480986 626614
rect 481542 626058 481574 626614
rect 480954 590614 481574 626058
rect 480954 590058 480986 590614
rect 481542 590058 481574 590614
rect 480954 554614 481574 590058
rect 480954 554058 480986 554614
rect 481542 554058 481574 554614
rect 480954 518614 481574 554058
rect 480954 518058 480986 518614
rect 481542 518058 481574 518614
rect 480954 482614 481574 518058
rect 480954 482058 480986 482614
rect 481542 482058 481574 482614
rect 480954 446614 481574 482058
rect 480954 446058 480986 446614
rect 481542 446058 481574 446614
rect 480954 410614 481574 446058
rect 480954 410058 480986 410614
rect 481542 410058 481574 410614
rect 480954 374614 481574 410058
rect 480954 374058 480986 374614
rect 481542 374058 481574 374614
rect 480954 338614 481574 374058
rect 480954 338058 480986 338614
rect 481542 338058 481574 338614
rect 480954 302614 481574 338058
rect 480954 302058 480986 302614
rect 481542 302058 481574 302614
rect 480954 266614 481574 302058
rect 480954 266058 480986 266614
rect 481542 266058 481574 266614
rect 480954 230614 481574 266058
rect 480954 230058 480986 230614
rect 481542 230058 481574 230614
rect 480954 194614 481574 230058
rect 480954 194058 480986 194614
rect 481542 194058 481574 194614
rect 480954 158614 481574 194058
rect 480954 158058 480986 158614
rect 481542 158058 481574 158614
rect 480954 122614 481574 158058
rect 480954 122058 480986 122614
rect 481542 122058 481574 122614
rect 480954 86614 481574 122058
rect 480954 86058 480986 86614
rect 481542 86058 481574 86614
rect 480954 50614 481574 86058
rect 480954 50058 480986 50614
rect 481542 50058 481574 50614
rect 480954 14614 481574 50058
rect 480954 14058 480986 14614
rect 481542 14058 481574 14614
rect 462954 -7622 462986 -7066
rect 463542 -7622 463574 -7066
rect 462954 -7654 463574 -7622
rect 480954 -6106 481574 14058
rect 487794 705798 488414 705830
rect 487794 705242 487826 705798
rect 488382 705242 488414 705798
rect 487794 669454 488414 705242
rect 487794 668898 487826 669454
rect 488382 668898 488414 669454
rect 487794 633454 488414 668898
rect 487794 632898 487826 633454
rect 488382 632898 488414 633454
rect 487794 597454 488414 632898
rect 487794 596898 487826 597454
rect 488382 596898 488414 597454
rect 487794 561454 488414 596898
rect 487794 560898 487826 561454
rect 488382 560898 488414 561454
rect 487794 525454 488414 560898
rect 487794 524898 487826 525454
rect 488382 524898 488414 525454
rect 487794 489454 488414 524898
rect 487794 488898 487826 489454
rect 488382 488898 488414 489454
rect 487794 453454 488414 488898
rect 487794 452898 487826 453454
rect 488382 452898 488414 453454
rect 487794 417454 488414 452898
rect 487794 416898 487826 417454
rect 488382 416898 488414 417454
rect 487794 381454 488414 416898
rect 487794 380898 487826 381454
rect 488382 380898 488414 381454
rect 487794 345454 488414 380898
rect 487794 344898 487826 345454
rect 488382 344898 488414 345454
rect 487794 309454 488414 344898
rect 487794 308898 487826 309454
rect 488382 308898 488414 309454
rect 487794 273454 488414 308898
rect 487794 272898 487826 273454
rect 488382 272898 488414 273454
rect 487794 237454 488414 272898
rect 487794 236898 487826 237454
rect 488382 236898 488414 237454
rect 487794 201454 488414 236898
rect 487794 200898 487826 201454
rect 488382 200898 488414 201454
rect 487794 165454 488414 200898
rect 487794 164898 487826 165454
rect 488382 164898 488414 165454
rect 487794 129454 488414 164898
rect 487794 128898 487826 129454
rect 488382 128898 488414 129454
rect 487794 93454 488414 128898
rect 487794 92898 487826 93454
rect 488382 92898 488414 93454
rect 487794 57454 488414 92898
rect 487794 56898 487826 57454
rect 488382 56898 488414 57454
rect 487794 21454 488414 56898
rect 487794 20898 487826 21454
rect 488382 20898 488414 21454
rect 487794 -1306 488414 20898
rect 487794 -1862 487826 -1306
rect 488382 -1862 488414 -1306
rect 487794 -1894 488414 -1862
rect 491514 673174 492134 707162
rect 491514 672618 491546 673174
rect 492102 672618 492134 673174
rect 491514 637174 492134 672618
rect 491514 636618 491546 637174
rect 492102 636618 492134 637174
rect 491514 601174 492134 636618
rect 491514 600618 491546 601174
rect 492102 600618 492134 601174
rect 491514 565174 492134 600618
rect 491514 564618 491546 565174
rect 492102 564618 492134 565174
rect 491514 529174 492134 564618
rect 491514 528618 491546 529174
rect 492102 528618 492134 529174
rect 491514 493174 492134 528618
rect 491514 492618 491546 493174
rect 492102 492618 492134 493174
rect 491514 457174 492134 492618
rect 491514 456618 491546 457174
rect 492102 456618 492134 457174
rect 491514 421174 492134 456618
rect 491514 420618 491546 421174
rect 492102 420618 492134 421174
rect 491514 385174 492134 420618
rect 491514 384618 491546 385174
rect 492102 384618 492134 385174
rect 491514 349174 492134 384618
rect 491514 348618 491546 349174
rect 492102 348618 492134 349174
rect 491514 313174 492134 348618
rect 491514 312618 491546 313174
rect 492102 312618 492134 313174
rect 491514 277174 492134 312618
rect 491514 276618 491546 277174
rect 492102 276618 492134 277174
rect 491514 241174 492134 276618
rect 491514 240618 491546 241174
rect 492102 240618 492134 241174
rect 491514 205174 492134 240618
rect 491514 204618 491546 205174
rect 492102 204618 492134 205174
rect 491514 169174 492134 204618
rect 491514 168618 491546 169174
rect 492102 168618 492134 169174
rect 491514 133174 492134 168618
rect 491514 132618 491546 133174
rect 492102 132618 492134 133174
rect 491514 97174 492134 132618
rect 491514 96618 491546 97174
rect 492102 96618 492134 97174
rect 491514 61174 492134 96618
rect 491514 60618 491546 61174
rect 492102 60618 492134 61174
rect 491514 25174 492134 60618
rect 491514 24618 491546 25174
rect 492102 24618 492134 25174
rect 491514 -3226 492134 24618
rect 491514 -3782 491546 -3226
rect 492102 -3782 492134 -3226
rect 491514 -3814 492134 -3782
rect 495234 676894 495854 709082
rect 495234 676338 495266 676894
rect 495822 676338 495854 676894
rect 495234 640894 495854 676338
rect 495234 640338 495266 640894
rect 495822 640338 495854 640894
rect 495234 604894 495854 640338
rect 495234 604338 495266 604894
rect 495822 604338 495854 604894
rect 495234 568894 495854 604338
rect 495234 568338 495266 568894
rect 495822 568338 495854 568894
rect 495234 532894 495854 568338
rect 495234 532338 495266 532894
rect 495822 532338 495854 532894
rect 495234 496894 495854 532338
rect 495234 496338 495266 496894
rect 495822 496338 495854 496894
rect 495234 460894 495854 496338
rect 495234 460338 495266 460894
rect 495822 460338 495854 460894
rect 495234 424894 495854 460338
rect 495234 424338 495266 424894
rect 495822 424338 495854 424894
rect 495234 388894 495854 424338
rect 495234 388338 495266 388894
rect 495822 388338 495854 388894
rect 495234 352894 495854 388338
rect 495234 352338 495266 352894
rect 495822 352338 495854 352894
rect 495234 316894 495854 352338
rect 495234 316338 495266 316894
rect 495822 316338 495854 316894
rect 495234 280894 495854 316338
rect 495234 280338 495266 280894
rect 495822 280338 495854 280894
rect 495234 244894 495854 280338
rect 495234 244338 495266 244894
rect 495822 244338 495854 244894
rect 495234 208894 495854 244338
rect 495234 208338 495266 208894
rect 495822 208338 495854 208894
rect 495234 172894 495854 208338
rect 495234 172338 495266 172894
rect 495822 172338 495854 172894
rect 495234 136894 495854 172338
rect 495234 136338 495266 136894
rect 495822 136338 495854 136894
rect 495234 100894 495854 136338
rect 495234 100338 495266 100894
rect 495822 100338 495854 100894
rect 495234 64894 495854 100338
rect 495234 64338 495266 64894
rect 495822 64338 495854 64894
rect 495234 28894 495854 64338
rect 495234 28338 495266 28894
rect 495822 28338 495854 28894
rect 495234 -5146 495854 28338
rect 495234 -5702 495266 -5146
rect 495822 -5702 495854 -5146
rect 495234 -5734 495854 -5702
rect 498954 680614 499574 711002
rect 516954 710598 517574 711590
rect 516954 710042 516986 710598
rect 517542 710042 517574 710598
rect 513234 708678 513854 709670
rect 513234 708122 513266 708678
rect 513822 708122 513854 708678
rect 509514 706758 510134 707750
rect 509514 706202 509546 706758
rect 510102 706202 510134 706758
rect 498954 680058 498986 680614
rect 499542 680058 499574 680614
rect 498954 644614 499574 680058
rect 498954 644058 498986 644614
rect 499542 644058 499574 644614
rect 498954 608614 499574 644058
rect 498954 608058 498986 608614
rect 499542 608058 499574 608614
rect 498954 572614 499574 608058
rect 498954 572058 498986 572614
rect 499542 572058 499574 572614
rect 498954 536614 499574 572058
rect 498954 536058 498986 536614
rect 499542 536058 499574 536614
rect 498954 500614 499574 536058
rect 498954 500058 498986 500614
rect 499542 500058 499574 500614
rect 498954 464614 499574 500058
rect 498954 464058 498986 464614
rect 499542 464058 499574 464614
rect 498954 428614 499574 464058
rect 498954 428058 498986 428614
rect 499542 428058 499574 428614
rect 498954 392614 499574 428058
rect 498954 392058 498986 392614
rect 499542 392058 499574 392614
rect 498954 356614 499574 392058
rect 498954 356058 498986 356614
rect 499542 356058 499574 356614
rect 498954 320614 499574 356058
rect 498954 320058 498986 320614
rect 499542 320058 499574 320614
rect 498954 284614 499574 320058
rect 498954 284058 498986 284614
rect 499542 284058 499574 284614
rect 498954 248614 499574 284058
rect 498954 248058 498986 248614
rect 499542 248058 499574 248614
rect 498954 212614 499574 248058
rect 498954 212058 498986 212614
rect 499542 212058 499574 212614
rect 498954 176614 499574 212058
rect 498954 176058 498986 176614
rect 499542 176058 499574 176614
rect 498954 140614 499574 176058
rect 498954 140058 498986 140614
rect 499542 140058 499574 140614
rect 498954 104614 499574 140058
rect 498954 104058 498986 104614
rect 499542 104058 499574 104614
rect 498954 68614 499574 104058
rect 498954 68058 498986 68614
rect 499542 68058 499574 68614
rect 498954 32614 499574 68058
rect 498954 32058 498986 32614
rect 499542 32058 499574 32614
rect 480954 -6662 480986 -6106
rect 481542 -6662 481574 -6106
rect 480954 -7654 481574 -6662
rect 498954 -7066 499574 32058
rect 505794 704838 506414 705830
rect 505794 704282 505826 704838
rect 506382 704282 506414 704838
rect 505794 687454 506414 704282
rect 505794 686898 505826 687454
rect 506382 686898 506414 687454
rect 505794 651454 506414 686898
rect 505794 650898 505826 651454
rect 506382 650898 506414 651454
rect 505794 615454 506414 650898
rect 505794 614898 505826 615454
rect 506382 614898 506414 615454
rect 505794 579454 506414 614898
rect 505794 578898 505826 579454
rect 506382 578898 506414 579454
rect 505794 543454 506414 578898
rect 505794 542898 505826 543454
rect 506382 542898 506414 543454
rect 505794 507454 506414 542898
rect 505794 506898 505826 507454
rect 506382 506898 506414 507454
rect 505794 471454 506414 506898
rect 505794 470898 505826 471454
rect 506382 470898 506414 471454
rect 505794 435454 506414 470898
rect 505794 434898 505826 435454
rect 506382 434898 506414 435454
rect 505794 399454 506414 434898
rect 505794 398898 505826 399454
rect 506382 398898 506414 399454
rect 505794 363454 506414 398898
rect 505794 362898 505826 363454
rect 506382 362898 506414 363454
rect 505794 327454 506414 362898
rect 505794 326898 505826 327454
rect 506382 326898 506414 327454
rect 505794 291454 506414 326898
rect 505794 290898 505826 291454
rect 506382 290898 506414 291454
rect 505794 255454 506414 290898
rect 505794 254898 505826 255454
rect 506382 254898 506414 255454
rect 505794 219454 506414 254898
rect 505794 218898 505826 219454
rect 506382 218898 506414 219454
rect 505794 183454 506414 218898
rect 505794 182898 505826 183454
rect 506382 182898 506414 183454
rect 505794 147454 506414 182898
rect 505794 146898 505826 147454
rect 506382 146898 506414 147454
rect 505794 111454 506414 146898
rect 505794 110898 505826 111454
rect 506382 110898 506414 111454
rect 505794 75454 506414 110898
rect 505794 74898 505826 75454
rect 506382 74898 506414 75454
rect 505794 39454 506414 74898
rect 505794 38898 505826 39454
rect 506382 38898 506414 39454
rect 505794 3454 506414 38898
rect 505794 2898 505826 3454
rect 506382 2898 506414 3454
rect 505794 -346 506414 2898
rect 505794 -902 505826 -346
rect 506382 -902 506414 -346
rect 505794 -1894 506414 -902
rect 509514 691174 510134 706202
rect 509514 690618 509546 691174
rect 510102 690618 510134 691174
rect 509514 655174 510134 690618
rect 509514 654618 509546 655174
rect 510102 654618 510134 655174
rect 509514 619174 510134 654618
rect 509514 618618 509546 619174
rect 510102 618618 510134 619174
rect 509514 583174 510134 618618
rect 509514 582618 509546 583174
rect 510102 582618 510134 583174
rect 509514 547174 510134 582618
rect 509514 546618 509546 547174
rect 510102 546618 510134 547174
rect 509514 511174 510134 546618
rect 509514 510618 509546 511174
rect 510102 510618 510134 511174
rect 509514 475174 510134 510618
rect 509514 474618 509546 475174
rect 510102 474618 510134 475174
rect 509514 439174 510134 474618
rect 509514 438618 509546 439174
rect 510102 438618 510134 439174
rect 509514 403174 510134 438618
rect 509514 402618 509546 403174
rect 510102 402618 510134 403174
rect 509514 367174 510134 402618
rect 509514 366618 509546 367174
rect 510102 366618 510134 367174
rect 509514 331174 510134 366618
rect 509514 330618 509546 331174
rect 510102 330618 510134 331174
rect 509514 295174 510134 330618
rect 509514 294618 509546 295174
rect 510102 294618 510134 295174
rect 509514 259174 510134 294618
rect 509514 258618 509546 259174
rect 510102 258618 510134 259174
rect 509514 223174 510134 258618
rect 509514 222618 509546 223174
rect 510102 222618 510134 223174
rect 509514 187174 510134 222618
rect 509514 186618 509546 187174
rect 510102 186618 510134 187174
rect 509514 151174 510134 186618
rect 509514 150618 509546 151174
rect 510102 150618 510134 151174
rect 509514 115174 510134 150618
rect 509514 114618 509546 115174
rect 510102 114618 510134 115174
rect 509514 79174 510134 114618
rect 509514 78618 509546 79174
rect 510102 78618 510134 79174
rect 509514 43174 510134 78618
rect 509514 42618 509546 43174
rect 510102 42618 510134 43174
rect 509514 7174 510134 42618
rect 509514 6618 509546 7174
rect 510102 6618 510134 7174
rect 509514 -2266 510134 6618
rect 509514 -2822 509546 -2266
rect 510102 -2822 510134 -2266
rect 509514 -3814 510134 -2822
rect 513234 694894 513854 708122
rect 513234 694338 513266 694894
rect 513822 694338 513854 694894
rect 513234 658894 513854 694338
rect 513234 658338 513266 658894
rect 513822 658338 513854 658894
rect 513234 622894 513854 658338
rect 513234 622338 513266 622894
rect 513822 622338 513854 622894
rect 513234 586894 513854 622338
rect 513234 586338 513266 586894
rect 513822 586338 513854 586894
rect 513234 550894 513854 586338
rect 513234 550338 513266 550894
rect 513822 550338 513854 550894
rect 513234 514894 513854 550338
rect 513234 514338 513266 514894
rect 513822 514338 513854 514894
rect 513234 478894 513854 514338
rect 513234 478338 513266 478894
rect 513822 478338 513854 478894
rect 513234 442894 513854 478338
rect 513234 442338 513266 442894
rect 513822 442338 513854 442894
rect 513234 406894 513854 442338
rect 513234 406338 513266 406894
rect 513822 406338 513854 406894
rect 513234 370894 513854 406338
rect 513234 370338 513266 370894
rect 513822 370338 513854 370894
rect 513234 334894 513854 370338
rect 513234 334338 513266 334894
rect 513822 334338 513854 334894
rect 513234 298894 513854 334338
rect 513234 298338 513266 298894
rect 513822 298338 513854 298894
rect 513234 262894 513854 298338
rect 513234 262338 513266 262894
rect 513822 262338 513854 262894
rect 513234 226894 513854 262338
rect 513234 226338 513266 226894
rect 513822 226338 513854 226894
rect 513234 190894 513854 226338
rect 513234 190338 513266 190894
rect 513822 190338 513854 190894
rect 513234 154894 513854 190338
rect 513234 154338 513266 154894
rect 513822 154338 513854 154894
rect 513234 118894 513854 154338
rect 513234 118338 513266 118894
rect 513822 118338 513854 118894
rect 513234 82894 513854 118338
rect 513234 82338 513266 82894
rect 513822 82338 513854 82894
rect 513234 46894 513854 82338
rect 513234 46338 513266 46894
rect 513822 46338 513854 46894
rect 513234 10894 513854 46338
rect 513234 10338 513266 10894
rect 513822 10338 513854 10894
rect 513234 -4186 513854 10338
rect 513234 -4742 513266 -4186
rect 513822 -4742 513854 -4186
rect 513234 -5734 513854 -4742
rect 516954 698614 517574 710042
rect 534954 711558 535574 711590
rect 534954 711002 534986 711558
rect 535542 711002 535574 711558
rect 531234 709638 531854 709670
rect 531234 709082 531266 709638
rect 531822 709082 531854 709638
rect 527514 707718 528134 707750
rect 527514 707162 527546 707718
rect 528102 707162 528134 707718
rect 516954 698058 516986 698614
rect 517542 698058 517574 698614
rect 516954 662614 517574 698058
rect 516954 662058 516986 662614
rect 517542 662058 517574 662614
rect 516954 626614 517574 662058
rect 516954 626058 516986 626614
rect 517542 626058 517574 626614
rect 516954 590614 517574 626058
rect 516954 590058 516986 590614
rect 517542 590058 517574 590614
rect 516954 554614 517574 590058
rect 516954 554058 516986 554614
rect 517542 554058 517574 554614
rect 516954 518614 517574 554058
rect 516954 518058 516986 518614
rect 517542 518058 517574 518614
rect 516954 482614 517574 518058
rect 516954 482058 516986 482614
rect 517542 482058 517574 482614
rect 516954 446614 517574 482058
rect 516954 446058 516986 446614
rect 517542 446058 517574 446614
rect 516954 410614 517574 446058
rect 516954 410058 516986 410614
rect 517542 410058 517574 410614
rect 516954 374614 517574 410058
rect 516954 374058 516986 374614
rect 517542 374058 517574 374614
rect 516954 338614 517574 374058
rect 516954 338058 516986 338614
rect 517542 338058 517574 338614
rect 516954 302614 517574 338058
rect 516954 302058 516986 302614
rect 517542 302058 517574 302614
rect 516954 266614 517574 302058
rect 516954 266058 516986 266614
rect 517542 266058 517574 266614
rect 516954 230614 517574 266058
rect 516954 230058 516986 230614
rect 517542 230058 517574 230614
rect 516954 194614 517574 230058
rect 516954 194058 516986 194614
rect 517542 194058 517574 194614
rect 516954 158614 517574 194058
rect 516954 158058 516986 158614
rect 517542 158058 517574 158614
rect 516954 122614 517574 158058
rect 516954 122058 516986 122614
rect 517542 122058 517574 122614
rect 516954 86614 517574 122058
rect 516954 86058 516986 86614
rect 517542 86058 517574 86614
rect 516954 50614 517574 86058
rect 516954 50058 516986 50614
rect 517542 50058 517574 50614
rect 516954 14614 517574 50058
rect 516954 14058 516986 14614
rect 517542 14058 517574 14614
rect 498954 -7622 498986 -7066
rect 499542 -7622 499574 -7066
rect 498954 -7654 499574 -7622
rect 516954 -6106 517574 14058
rect 523794 705798 524414 705830
rect 523794 705242 523826 705798
rect 524382 705242 524414 705798
rect 523794 669454 524414 705242
rect 523794 668898 523826 669454
rect 524382 668898 524414 669454
rect 523794 633454 524414 668898
rect 523794 632898 523826 633454
rect 524382 632898 524414 633454
rect 523794 597454 524414 632898
rect 523794 596898 523826 597454
rect 524382 596898 524414 597454
rect 523794 561454 524414 596898
rect 523794 560898 523826 561454
rect 524382 560898 524414 561454
rect 523794 525454 524414 560898
rect 523794 524898 523826 525454
rect 524382 524898 524414 525454
rect 523794 489454 524414 524898
rect 523794 488898 523826 489454
rect 524382 488898 524414 489454
rect 523794 453454 524414 488898
rect 523794 452898 523826 453454
rect 524382 452898 524414 453454
rect 523794 417454 524414 452898
rect 523794 416898 523826 417454
rect 524382 416898 524414 417454
rect 523794 381454 524414 416898
rect 523794 380898 523826 381454
rect 524382 380898 524414 381454
rect 523794 345454 524414 380898
rect 523794 344898 523826 345454
rect 524382 344898 524414 345454
rect 523794 309454 524414 344898
rect 523794 308898 523826 309454
rect 524382 308898 524414 309454
rect 523794 273454 524414 308898
rect 523794 272898 523826 273454
rect 524382 272898 524414 273454
rect 523794 237454 524414 272898
rect 523794 236898 523826 237454
rect 524382 236898 524414 237454
rect 523794 201454 524414 236898
rect 523794 200898 523826 201454
rect 524382 200898 524414 201454
rect 523794 165454 524414 200898
rect 523794 164898 523826 165454
rect 524382 164898 524414 165454
rect 523794 129454 524414 164898
rect 523794 128898 523826 129454
rect 524382 128898 524414 129454
rect 523794 93454 524414 128898
rect 523794 92898 523826 93454
rect 524382 92898 524414 93454
rect 523794 57454 524414 92898
rect 523794 56898 523826 57454
rect 524382 56898 524414 57454
rect 523794 21454 524414 56898
rect 523794 20898 523826 21454
rect 524382 20898 524414 21454
rect 523794 -1306 524414 20898
rect 523794 -1862 523826 -1306
rect 524382 -1862 524414 -1306
rect 523794 -1894 524414 -1862
rect 527514 673174 528134 707162
rect 527514 672618 527546 673174
rect 528102 672618 528134 673174
rect 527514 637174 528134 672618
rect 527514 636618 527546 637174
rect 528102 636618 528134 637174
rect 527514 601174 528134 636618
rect 527514 600618 527546 601174
rect 528102 600618 528134 601174
rect 527514 565174 528134 600618
rect 527514 564618 527546 565174
rect 528102 564618 528134 565174
rect 527514 529174 528134 564618
rect 527514 528618 527546 529174
rect 528102 528618 528134 529174
rect 527514 493174 528134 528618
rect 527514 492618 527546 493174
rect 528102 492618 528134 493174
rect 527514 457174 528134 492618
rect 527514 456618 527546 457174
rect 528102 456618 528134 457174
rect 527514 421174 528134 456618
rect 527514 420618 527546 421174
rect 528102 420618 528134 421174
rect 527514 385174 528134 420618
rect 527514 384618 527546 385174
rect 528102 384618 528134 385174
rect 527514 349174 528134 384618
rect 527514 348618 527546 349174
rect 528102 348618 528134 349174
rect 527514 313174 528134 348618
rect 527514 312618 527546 313174
rect 528102 312618 528134 313174
rect 527514 277174 528134 312618
rect 527514 276618 527546 277174
rect 528102 276618 528134 277174
rect 527514 241174 528134 276618
rect 527514 240618 527546 241174
rect 528102 240618 528134 241174
rect 527514 205174 528134 240618
rect 527514 204618 527546 205174
rect 528102 204618 528134 205174
rect 527514 169174 528134 204618
rect 527514 168618 527546 169174
rect 528102 168618 528134 169174
rect 527514 133174 528134 168618
rect 527514 132618 527546 133174
rect 528102 132618 528134 133174
rect 527514 97174 528134 132618
rect 527514 96618 527546 97174
rect 528102 96618 528134 97174
rect 527514 61174 528134 96618
rect 527514 60618 527546 61174
rect 528102 60618 528134 61174
rect 527514 25174 528134 60618
rect 527514 24618 527546 25174
rect 528102 24618 528134 25174
rect 527514 -3226 528134 24618
rect 527514 -3782 527546 -3226
rect 528102 -3782 528134 -3226
rect 527514 -3814 528134 -3782
rect 531234 676894 531854 709082
rect 531234 676338 531266 676894
rect 531822 676338 531854 676894
rect 531234 640894 531854 676338
rect 531234 640338 531266 640894
rect 531822 640338 531854 640894
rect 531234 604894 531854 640338
rect 531234 604338 531266 604894
rect 531822 604338 531854 604894
rect 531234 568894 531854 604338
rect 531234 568338 531266 568894
rect 531822 568338 531854 568894
rect 531234 532894 531854 568338
rect 531234 532338 531266 532894
rect 531822 532338 531854 532894
rect 531234 496894 531854 532338
rect 531234 496338 531266 496894
rect 531822 496338 531854 496894
rect 531234 460894 531854 496338
rect 531234 460338 531266 460894
rect 531822 460338 531854 460894
rect 531234 424894 531854 460338
rect 531234 424338 531266 424894
rect 531822 424338 531854 424894
rect 531234 388894 531854 424338
rect 531234 388338 531266 388894
rect 531822 388338 531854 388894
rect 531234 352894 531854 388338
rect 531234 352338 531266 352894
rect 531822 352338 531854 352894
rect 531234 316894 531854 352338
rect 531234 316338 531266 316894
rect 531822 316338 531854 316894
rect 531234 280894 531854 316338
rect 531234 280338 531266 280894
rect 531822 280338 531854 280894
rect 531234 244894 531854 280338
rect 531234 244338 531266 244894
rect 531822 244338 531854 244894
rect 531234 208894 531854 244338
rect 531234 208338 531266 208894
rect 531822 208338 531854 208894
rect 531234 172894 531854 208338
rect 531234 172338 531266 172894
rect 531822 172338 531854 172894
rect 531234 136894 531854 172338
rect 531234 136338 531266 136894
rect 531822 136338 531854 136894
rect 531234 100894 531854 136338
rect 531234 100338 531266 100894
rect 531822 100338 531854 100894
rect 531234 64894 531854 100338
rect 531234 64338 531266 64894
rect 531822 64338 531854 64894
rect 531234 28894 531854 64338
rect 531234 28338 531266 28894
rect 531822 28338 531854 28894
rect 531234 -5146 531854 28338
rect 531234 -5702 531266 -5146
rect 531822 -5702 531854 -5146
rect 531234 -5734 531854 -5702
rect 534954 680614 535574 711002
rect 552954 710598 553574 711590
rect 552954 710042 552986 710598
rect 553542 710042 553574 710598
rect 549234 708678 549854 709670
rect 549234 708122 549266 708678
rect 549822 708122 549854 708678
rect 545514 706758 546134 707750
rect 545514 706202 545546 706758
rect 546102 706202 546134 706758
rect 534954 680058 534986 680614
rect 535542 680058 535574 680614
rect 534954 644614 535574 680058
rect 534954 644058 534986 644614
rect 535542 644058 535574 644614
rect 534954 608614 535574 644058
rect 534954 608058 534986 608614
rect 535542 608058 535574 608614
rect 534954 572614 535574 608058
rect 534954 572058 534986 572614
rect 535542 572058 535574 572614
rect 534954 536614 535574 572058
rect 534954 536058 534986 536614
rect 535542 536058 535574 536614
rect 534954 500614 535574 536058
rect 534954 500058 534986 500614
rect 535542 500058 535574 500614
rect 534954 464614 535574 500058
rect 534954 464058 534986 464614
rect 535542 464058 535574 464614
rect 534954 428614 535574 464058
rect 534954 428058 534986 428614
rect 535542 428058 535574 428614
rect 534954 392614 535574 428058
rect 534954 392058 534986 392614
rect 535542 392058 535574 392614
rect 534954 356614 535574 392058
rect 534954 356058 534986 356614
rect 535542 356058 535574 356614
rect 534954 320614 535574 356058
rect 534954 320058 534986 320614
rect 535542 320058 535574 320614
rect 534954 284614 535574 320058
rect 534954 284058 534986 284614
rect 535542 284058 535574 284614
rect 534954 248614 535574 284058
rect 534954 248058 534986 248614
rect 535542 248058 535574 248614
rect 534954 212614 535574 248058
rect 534954 212058 534986 212614
rect 535542 212058 535574 212614
rect 534954 176614 535574 212058
rect 534954 176058 534986 176614
rect 535542 176058 535574 176614
rect 534954 140614 535574 176058
rect 534954 140058 534986 140614
rect 535542 140058 535574 140614
rect 534954 104614 535574 140058
rect 534954 104058 534986 104614
rect 535542 104058 535574 104614
rect 534954 68614 535574 104058
rect 534954 68058 534986 68614
rect 535542 68058 535574 68614
rect 534954 32614 535574 68058
rect 534954 32058 534986 32614
rect 535542 32058 535574 32614
rect 516954 -6662 516986 -6106
rect 517542 -6662 517574 -6106
rect 516954 -7654 517574 -6662
rect 534954 -7066 535574 32058
rect 541794 704838 542414 705830
rect 541794 704282 541826 704838
rect 542382 704282 542414 704838
rect 541794 687454 542414 704282
rect 541794 686898 541826 687454
rect 542382 686898 542414 687454
rect 541794 651454 542414 686898
rect 541794 650898 541826 651454
rect 542382 650898 542414 651454
rect 541794 615454 542414 650898
rect 541794 614898 541826 615454
rect 542382 614898 542414 615454
rect 541794 579454 542414 614898
rect 541794 578898 541826 579454
rect 542382 578898 542414 579454
rect 541794 543454 542414 578898
rect 541794 542898 541826 543454
rect 542382 542898 542414 543454
rect 541794 507454 542414 542898
rect 541794 506898 541826 507454
rect 542382 506898 542414 507454
rect 541794 471454 542414 506898
rect 541794 470898 541826 471454
rect 542382 470898 542414 471454
rect 541794 435454 542414 470898
rect 541794 434898 541826 435454
rect 542382 434898 542414 435454
rect 541794 399454 542414 434898
rect 541794 398898 541826 399454
rect 542382 398898 542414 399454
rect 541794 363454 542414 398898
rect 541794 362898 541826 363454
rect 542382 362898 542414 363454
rect 541794 327454 542414 362898
rect 541794 326898 541826 327454
rect 542382 326898 542414 327454
rect 541794 291454 542414 326898
rect 541794 290898 541826 291454
rect 542382 290898 542414 291454
rect 541794 255454 542414 290898
rect 541794 254898 541826 255454
rect 542382 254898 542414 255454
rect 541794 219454 542414 254898
rect 541794 218898 541826 219454
rect 542382 218898 542414 219454
rect 541794 183454 542414 218898
rect 541794 182898 541826 183454
rect 542382 182898 542414 183454
rect 541794 147454 542414 182898
rect 541794 146898 541826 147454
rect 542382 146898 542414 147454
rect 541794 111454 542414 146898
rect 541794 110898 541826 111454
rect 542382 110898 542414 111454
rect 541794 75454 542414 110898
rect 541794 74898 541826 75454
rect 542382 74898 542414 75454
rect 541794 39454 542414 74898
rect 541794 38898 541826 39454
rect 542382 38898 542414 39454
rect 541794 3454 542414 38898
rect 541794 2898 541826 3454
rect 542382 2898 542414 3454
rect 541794 -346 542414 2898
rect 541794 -902 541826 -346
rect 542382 -902 542414 -346
rect 541794 -1894 542414 -902
rect 545514 691174 546134 706202
rect 545514 690618 545546 691174
rect 546102 690618 546134 691174
rect 545514 655174 546134 690618
rect 545514 654618 545546 655174
rect 546102 654618 546134 655174
rect 545514 619174 546134 654618
rect 545514 618618 545546 619174
rect 546102 618618 546134 619174
rect 545514 583174 546134 618618
rect 545514 582618 545546 583174
rect 546102 582618 546134 583174
rect 545514 547174 546134 582618
rect 545514 546618 545546 547174
rect 546102 546618 546134 547174
rect 545514 511174 546134 546618
rect 545514 510618 545546 511174
rect 546102 510618 546134 511174
rect 545514 475174 546134 510618
rect 545514 474618 545546 475174
rect 546102 474618 546134 475174
rect 545514 439174 546134 474618
rect 545514 438618 545546 439174
rect 546102 438618 546134 439174
rect 545514 403174 546134 438618
rect 545514 402618 545546 403174
rect 546102 402618 546134 403174
rect 545514 367174 546134 402618
rect 545514 366618 545546 367174
rect 546102 366618 546134 367174
rect 545514 331174 546134 366618
rect 545514 330618 545546 331174
rect 546102 330618 546134 331174
rect 545514 295174 546134 330618
rect 545514 294618 545546 295174
rect 546102 294618 546134 295174
rect 545514 259174 546134 294618
rect 545514 258618 545546 259174
rect 546102 258618 546134 259174
rect 545514 223174 546134 258618
rect 545514 222618 545546 223174
rect 546102 222618 546134 223174
rect 545514 187174 546134 222618
rect 545514 186618 545546 187174
rect 546102 186618 546134 187174
rect 545514 151174 546134 186618
rect 545514 150618 545546 151174
rect 546102 150618 546134 151174
rect 545514 115174 546134 150618
rect 545514 114618 545546 115174
rect 546102 114618 546134 115174
rect 545514 79174 546134 114618
rect 545514 78618 545546 79174
rect 546102 78618 546134 79174
rect 545514 43174 546134 78618
rect 545514 42618 545546 43174
rect 546102 42618 546134 43174
rect 545514 7174 546134 42618
rect 545514 6618 545546 7174
rect 546102 6618 546134 7174
rect 545514 -2266 546134 6618
rect 545514 -2822 545546 -2266
rect 546102 -2822 546134 -2266
rect 545514 -3814 546134 -2822
rect 549234 694894 549854 708122
rect 549234 694338 549266 694894
rect 549822 694338 549854 694894
rect 549234 658894 549854 694338
rect 549234 658338 549266 658894
rect 549822 658338 549854 658894
rect 549234 622894 549854 658338
rect 549234 622338 549266 622894
rect 549822 622338 549854 622894
rect 549234 586894 549854 622338
rect 549234 586338 549266 586894
rect 549822 586338 549854 586894
rect 549234 550894 549854 586338
rect 549234 550338 549266 550894
rect 549822 550338 549854 550894
rect 549234 514894 549854 550338
rect 549234 514338 549266 514894
rect 549822 514338 549854 514894
rect 549234 478894 549854 514338
rect 549234 478338 549266 478894
rect 549822 478338 549854 478894
rect 549234 442894 549854 478338
rect 549234 442338 549266 442894
rect 549822 442338 549854 442894
rect 549234 406894 549854 442338
rect 549234 406338 549266 406894
rect 549822 406338 549854 406894
rect 549234 370894 549854 406338
rect 549234 370338 549266 370894
rect 549822 370338 549854 370894
rect 549234 334894 549854 370338
rect 549234 334338 549266 334894
rect 549822 334338 549854 334894
rect 549234 298894 549854 334338
rect 549234 298338 549266 298894
rect 549822 298338 549854 298894
rect 549234 262894 549854 298338
rect 549234 262338 549266 262894
rect 549822 262338 549854 262894
rect 549234 226894 549854 262338
rect 549234 226338 549266 226894
rect 549822 226338 549854 226894
rect 549234 190894 549854 226338
rect 549234 190338 549266 190894
rect 549822 190338 549854 190894
rect 549234 154894 549854 190338
rect 549234 154338 549266 154894
rect 549822 154338 549854 154894
rect 549234 118894 549854 154338
rect 549234 118338 549266 118894
rect 549822 118338 549854 118894
rect 549234 82894 549854 118338
rect 549234 82338 549266 82894
rect 549822 82338 549854 82894
rect 549234 46894 549854 82338
rect 549234 46338 549266 46894
rect 549822 46338 549854 46894
rect 549234 10894 549854 46338
rect 549234 10338 549266 10894
rect 549822 10338 549854 10894
rect 549234 -4186 549854 10338
rect 549234 -4742 549266 -4186
rect 549822 -4742 549854 -4186
rect 549234 -5734 549854 -4742
rect 552954 698614 553574 710042
rect 570954 711558 571574 711590
rect 570954 711002 570986 711558
rect 571542 711002 571574 711558
rect 567234 709638 567854 709670
rect 567234 709082 567266 709638
rect 567822 709082 567854 709638
rect 563514 707718 564134 707750
rect 563514 707162 563546 707718
rect 564102 707162 564134 707718
rect 552954 698058 552986 698614
rect 553542 698058 553574 698614
rect 552954 662614 553574 698058
rect 552954 662058 552986 662614
rect 553542 662058 553574 662614
rect 552954 626614 553574 662058
rect 552954 626058 552986 626614
rect 553542 626058 553574 626614
rect 552954 590614 553574 626058
rect 552954 590058 552986 590614
rect 553542 590058 553574 590614
rect 552954 554614 553574 590058
rect 552954 554058 552986 554614
rect 553542 554058 553574 554614
rect 552954 518614 553574 554058
rect 552954 518058 552986 518614
rect 553542 518058 553574 518614
rect 552954 482614 553574 518058
rect 552954 482058 552986 482614
rect 553542 482058 553574 482614
rect 552954 446614 553574 482058
rect 552954 446058 552986 446614
rect 553542 446058 553574 446614
rect 552954 410614 553574 446058
rect 552954 410058 552986 410614
rect 553542 410058 553574 410614
rect 552954 374614 553574 410058
rect 552954 374058 552986 374614
rect 553542 374058 553574 374614
rect 552954 338614 553574 374058
rect 552954 338058 552986 338614
rect 553542 338058 553574 338614
rect 552954 302614 553574 338058
rect 552954 302058 552986 302614
rect 553542 302058 553574 302614
rect 552954 266614 553574 302058
rect 552954 266058 552986 266614
rect 553542 266058 553574 266614
rect 552954 230614 553574 266058
rect 552954 230058 552986 230614
rect 553542 230058 553574 230614
rect 552954 194614 553574 230058
rect 552954 194058 552986 194614
rect 553542 194058 553574 194614
rect 552954 158614 553574 194058
rect 552954 158058 552986 158614
rect 553542 158058 553574 158614
rect 552954 122614 553574 158058
rect 552954 122058 552986 122614
rect 553542 122058 553574 122614
rect 552954 86614 553574 122058
rect 552954 86058 552986 86614
rect 553542 86058 553574 86614
rect 552954 50614 553574 86058
rect 552954 50058 552986 50614
rect 553542 50058 553574 50614
rect 552954 14614 553574 50058
rect 552954 14058 552986 14614
rect 553542 14058 553574 14614
rect 534954 -7622 534986 -7066
rect 535542 -7622 535574 -7066
rect 534954 -7654 535574 -7622
rect 552954 -6106 553574 14058
rect 559794 705798 560414 705830
rect 559794 705242 559826 705798
rect 560382 705242 560414 705798
rect 559794 669454 560414 705242
rect 559794 668898 559826 669454
rect 560382 668898 560414 669454
rect 559794 633454 560414 668898
rect 559794 632898 559826 633454
rect 560382 632898 560414 633454
rect 559794 597454 560414 632898
rect 559794 596898 559826 597454
rect 560382 596898 560414 597454
rect 559794 561454 560414 596898
rect 559794 560898 559826 561454
rect 560382 560898 560414 561454
rect 559794 525454 560414 560898
rect 559794 524898 559826 525454
rect 560382 524898 560414 525454
rect 559794 489454 560414 524898
rect 559794 488898 559826 489454
rect 560382 488898 560414 489454
rect 559794 453454 560414 488898
rect 559794 452898 559826 453454
rect 560382 452898 560414 453454
rect 559794 417454 560414 452898
rect 559794 416898 559826 417454
rect 560382 416898 560414 417454
rect 559794 381454 560414 416898
rect 559794 380898 559826 381454
rect 560382 380898 560414 381454
rect 559794 345454 560414 380898
rect 559794 344898 559826 345454
rect 560382 344898 560414 345454
rect 559794 309454 560414 344898
rect 559794 308898 559826 309454
rect 560382 308898 560414 309454
rect 559794 273454 560414 308898
rect 559794 272898 559826 273454
rect 560382 272898 560414 273454
rect 559794 237454 560414 272898
rect 559794 236898 559826 237454
rect 560382 236898 560414 237454
rect 559794 201454 560414 236898
rect 559794 200898 559826 201454
rect 560382 200898 560414 201454
rect 559794 165454 560414 200898
rect 559794 164898 559826 165454
rect 560382 164898 560414 165454
rect 559794 129454 560414 164898
rect 559794 128898 559826 129454
rect 560382 128898 560414 129454
rect 559794 93454 560414 128898
rect 559794 92898 559826 93454
rect 560382 92898 560414 93454
rect 559794 57454 560414 92898
rect 559794 56898 559826 57454
rect 560382 56898 560414 57454
rect 559794 21454 560414 56898
rect 559794 20898 559826 21454
rect 560382 20898 560414 21454
rect 559794 -1306 560414 20898
rect 559794 -1862 559826 -1306
rect 560382 -1862 560414 -1306
rect 559794 -1894 560414 -1862
rect 563514 673174 564134 707162
rect 563514 672618 563546 673174
rect 564102 672618 564134 673174
rect 563514 637174 564134 672618
rect 563514 636618 563546 637174
rect 564102 636618 564134 637174
rect 563514 601174 564134 636618
rect 563514 600618 563546 601174
rect 564102 600618 564134 601174
rect 563514 565174 564134 600618
rect 563514 564618 563546 565174
rect 564102 564618 564134 565174
rect 563514 529174 564134 564618
rect 563514 528618 563546 529174
rect 564102 528618 564134 529174
rect 563514 493174 564134 528618
rect 563514 492618 563546 493174
rect 564102 492618 564134 493174
rect 563514 457174 564134 492618
rect 563514 456618 563546 457174
rect 564102 456618 564134 457174
rect 563514 421174 564134 456618
rect 563514 420618 563546 421174
rect 564102 420618 564134 421174
rect 563514 385174 564134 420618
rect 563514 384618 563546 385174
rect 564102 384618 564134 385174
rect 563514 349174 564134 384618
rect 563514 348618 563546 349174
rect 564102 348618 564134 349174
rect 563514 313174 564134 348618
rect 563514 312618 563546 313174
rect 564102 312618 564134 313174
rect 563514 277174 564134 312618
rect 563514 276618 563546 277174
rect 564102 276618 564134 277174
rect 563514 241174 564134 276618
rect 563514 240618 563546 241174
rect 564102 240618 564134 241174
rect 563514 205174 564134 240618
rect 563514 204618 563546 205174
rect 564102 204618 564134 205174
rect 563514 169174 564134 204618
rect 563514 168618 563546 169174
rect 564102 168618 564134 169174
rect 563514 133174 564134 168618
rect 563514 132618 563546 133174
rect 564102 132618 564134 133174
rect 563514 97174 564134 132618
rect 563514 96618 563546 97174
rect 564102 96618 564134 97174
rect 563514 61174 564134 96618
rect 563514 60618 563546 61174
rect 564102 60618 564134 61174
rect 563514 25174 564134 60618
rect 563514 24618 563546 25174
rect 564102 24618 564134 25174
rect 563514 -3226 564134 24618
rect 563514 -3782 563546 -3226
rect 564102 -3782 564134 -3226
rect 563514 -3814 564134 -3782
rect 567234 676894 567854 709082
rect 567234 676338 567266 676894
rect 567822 676338 567854 676894
rect 567234 640894 567854 676338
rect 567234 640338 567266 640894
rect 567822 640338 567854 640894
rect 567234 604894 567854 640338
rect 567234 604338 567266 604894
rect 567822 604338 567854 604894
rect 567234 568894 567854 604338
rect 567234 568338 567266 568894
rect 567822 568338 567854 568894
rect 567234 532894 567854 568338
rect 567234 532338 567266 532894
rect 567822 532338 567854 532894
rect 567234 496894 567854 532338
rect 567234 496338 567266 496894
rect 567822 496338 567854 496894
rect 567234 460894 567854 496338
rect 567234 460338 567266 460894
rect 567822 460338 567854 460894
rect 567234 424894 567854 460338
rect 567234 424338 567266 424894
rect 567822 424338 567854 424894
rect 567234 388894 567854 424338
rect 567234 388338 567266 388894
rect 567822 388338 567854 388894
rect 567234 352894 567854 388338
rect 567234 352338 567266 352894
rect 567822 352338 567854 352894
rect 567234 316894 567854 352338
rect 567234 316338 567266 316894
rect 567822 316338 567854 316894
rect 567234 280894 567854 316338
rect 567234 280338 567266 280894
rect 567822 280338 567854 280894
rect 567234 244894 567854 280338
rect 567234 244338 567266 244894
rect 567822 244338 567854 244894
rect 567234 208894 567854 244338
rect 567234 208338 567266 208894
rect 567822 208338 567854 208894
rect 567234 172894 567854 208338
rect 567234 172338 567266 172894
rect 567822 172338 567854 172894
rect 567234 136894 567854 172338
rect 567234 136338 567266 136894
rect 567822 136338 567854 136894
rect 567234 100894 567854 136338
rect 567234 100338 567266 100894
rect 567822 100338 567854 100894
rect 567234 64894 567854 100338
rect 567234 64338 567266 64894
rect 567822 64338 567854 64894
rect 567234 28894 567854 64338
rect 567234 28338 567266 28894
rect 567822 28338 567854 28894
rect 567234 -5146 567854 28338
rect 567234 -5702 567266 -5146
rect 567822 -5702 567854 -5146
rect 567234 -5734 567854 -5702
rect 570954 680614 571574 711002
rect 592030 711558 592650 711590
rect 592030 711002 592062 711558
rect 592618 711002 592650 711558
rect 591070 710598 591690 710630
rect 591070 710042 591102 710598
rect 591658 710042 591690 710598
rect 590110 709638 590730 709670
rect 590110 709082 590142 709638
rect 590698 709082 590730 709638
rect 589150 708678 589770 708710
rect 589150 708122 589182 708678
rect 589738 708122 589770 708678
rect 581514 706758 582134 707750
rect 588190 707718 588810 707750
rect 588190 707162 588222 707718
rect 588778 707162 588810 707718
rect 581514 706202 581546 706758
rect 582102 706202 582134 706758
rect 570954 680058 570986 680614
rect 571542 680058 571574 680614
rect 570954 644614 571574 680058
rect 570954 644058 570986 644614
rect 571542 644058 571574 644614
rect 570954 608614 571574 644058
rect 570954 608058 570986 608614
rect 571542 608058 571574 608614
rect 570954 572614 571574 608058
rect 570954 572058 570986 572614
rect 571542 572058 571574 572614
rect 570954 536614 571574 572058
rect 570954 536058 570986 536614
rect 571542 536058 571574 536614
rect 570954 500614 571574 536058
rect 570954 500058 570986 500614
rect 571542 500058 571574 500614
rect 570954 464614 571574 500058
rect 570954 464058 570986 464614
rect 571542 464058 571574 464614
rect 570954 428614 571574 464058
rect 570954 428058 570986 428614
rect 571542 428058 571574 428614
rect 570954 392614 571574 428058
rect 570954 392058 570986 392614
rect 571542 392058 571574 392614
rect 570954 356614 571574 392058
rect 570954 356058 570986 356614
rect 571542 356058 571574 356614
rect 570954 320614 571574 356058
rect 570954 320058 570986 320614
rect 571542 320058 571574 320614
rect 570954 284614 571574 320058
rect 570954 284058 570986 284614
rect 571542 284058 571574 284614
rect 570954 248614 571574 284058
rect 570954 248058 570986 248614
rect 571542 248058 571574 248614
rect 570954 212614 571574 248058
rect 570954 212058 570986 212614
rect 571542 212058 571574 212614
rect 570954 176614 571574 212058
rect 570954 176058 570986 176614
rect 571542 176058 571574 176614
rect 570954 140614 571574 176058
rect 570954 140058 570986 140614
rect 571542 140058 571574 140614
rect 570954 104614 571574 140058
rect 570954 104058 570986 104614
rect 571542 104058 571574 104614
rect 570954 68614 571574 104058
rect 570954 68058 570986 68614
rect 571542 68058 571574 68614
rect 570954 32614 571574 68058
rect 570954 32058 570986 32614
rect 571542 32058 571574 32614
rect 552954 -6662 552986 -6106
rect 553542 -6662 553574 -6106
rect 552954 -7654 553574 -6662
rect 570954 -7066 571574 32058
rect 577794 704838 578414 705830
rect 577794 704282 577826 704838
rect 578382 704282 578414 704838
rect 577794 687454 578414 704282
rect 577794 686898 577826 687454
rect 578382 686898 578414 687454
rect 577794 651454 578414 686898
rect 577794 650898 577826 651454
rect 578382 650898 578414 651454
rect 577794 615454 578414 650898
rect 577794 614898 577826 615454
rect 578382 614898 578414 615454
rect 577794 579454 578414 614898
rect 577794 578898 577826 579454
rect 578382 578898 578414 579454
rect 577794 543454 578414 578898
rect 577794 542898 577826 543454
rect 578382 542898 578414 543454
rect 577794 507454 578414 542898
rect 577794 506898 577826 507454
rect 578382 506898 578414 507454
rect 577794 471454 578414 506898
rect 577794 470898 577826 471454
rect 578382 470898 578414 471454
rect 577794 435454 578414 470898
rect 577794 434898 577826 435454
rect 578382 434898 578414 435454
rect 577794 399454 578414 434898
rect 577794 398898 577826 399454
rect 578382 398898 578414 399454
rect 577794 363454 578414 398898
rect 577794 362898 577826 363454
rect 578382 362898 578414 363454
rect 577794 327454 578414 362898
rect 577794 326898 577826 327454
rect 578382 326898 578414 327454
rect 577794 291454 578414 326898
rect 577794 290898 577826 291454
rect 578382 290898 578414 291454
rect 577794 255454 578414 290898
rect 577794 254898 577826 255454
rect 578382 254898 578414 255454
rect 577794 219454 578414 254898
rect 577794 218898 577826 219454
rect 578382 218898 578414 219454
rect 577794 183454 578414 218898
rect 577794 182898 577826 183454
rect 578382 182898 578414 183454
rect 577794 147454 578414 182898
rect 577794 146898 577826 147454
rect 578382 146898 578414 147454
rect 577794 111454 578414 146898
rect 577794 110898 577826 111454
rect 578382 110898 578414 111454
rect 577794 75454 578414 110898
rect 577794 74898 577826 75454
rect 578382 74898 578414 75454
rect 577794 39454 578414 74898
rect 577794 38898 577826 39454
rect 578382 38898 578414 39454
rect 577794 3454 578414 38898
rect 577794 2898 577826 3454
rect 578382 2898 578414 3454
rect 577794 -346 578414 2898
rect 577794 -902 577826 -346
rect 578382 -902 578414 -346
rect 577794 -1894 578414 -902
rect 581514 691174 582134 706202
rect 587230 706758 587850 706790
rect 587230 706202 587262 706758
rect 587818 706202 587850 706758
rect 586270 705798 586890 705830
rect 586270 705242 586302 705798
rect 586858 705242 586890 705798
rect 581514 690618 581546 691174
rect 582102 690618 582134 691174
rect 581514 655174 582134 690618
rect 581514 654618 581546 655174
rect 582102 654618 582134 655174
rect 581514 619174 582134 654618
rect 581514 618618 581546 619174
rect 582102 618618 582134 619174
rect 581514 583174 582134 618618
rect 581514 582618 581546 583174
rect 582102 582618 582134 583174
rect 581514 547174 582134 582618
rect 581514 546618 581546 547174
rect 582102 546618 582134 547174
rect 581514 511174 582134 546618
rect 581514 510618 581546 511174
rect 582102 510618 582134 511174
rect 581514 475174 582134 510618
rect 581514 474618 581546 475174
rect 582102 474618 582134 475174
rect 581514 439174 582134 474618
rect 581514 438618 581546 439174
rect 582102 438618 582134 439174
rect 581514 403174 582134 438618
rect 581514 402618 581546 403174
rect 582102 402618 582134 403174
rect 581514 367174 582134 402618
rect 581514 366618 581546 367174
rect 582102 366618 582134 367174
rect 581514 331174 582134 366618
rect 581514 330618 581546 331174
rect 582102 330618 582134 331174
rect 581514 295174 582134 330618
rect 581514 294618 581546 295174
rect 582102 294618 582134 295174
rect 581514 259174 582134 294618
rect 581514 258618 581546 259174
rect 582102 258618 582134 259174
rect 581514 223174 582134 258618
rect 581514 222618 581546 223174
rect 582102 222618 582134 223174
rect 581514 187174 582134 222618
rect 581514 186618 581546 187174
rect 582102 186618 582134 187174
rect 581514 151174 582134 186618
rect 581514 150618 581546 151174
rect 582102 150618 582134 151174
rect 581514 115174 582134 150618
rect 581514 114618 581546 115174
rect 582102 114618 582134 115174
rect 581514 79174 582134 114618
rect 581514 78618 581546 79174
rect 582102 78618 582134 79174
rect 581514 43174 582134 78618
rect 581514 42618 581546 43174
rect 582102 42618 582134 43174
rect 581514 7174 582134 42618
rect 581514 6618 581546 7174
rect 582102 6618 582134 7174
rect 581514 -2266 582134 6618
rect 585310 704838 585930 704870
rect 585310 704282 585342 704838
rect 585898 704282 585930 704838
rect 585310 687454 585930 704282
rect 585310 686898 585342 687454
rect 585898 686898 585930 687454
rect 585310 651454 585930 686898
rect 585310 650898 585342 651454
rect 585898 650898 585930 651454
rect 585310 615454 585930 650898
rect 585310 614898 585342 615454
rect 585898 614898 585930 615454
rect 585310 579454 585930 614898
rect 585310 578898 585342 579454
rect 585898 578898 585930 579454
rect 585310 543454 585930 578898
rect 585310 542898 585342 543454
rect 585898 542898 585930 543454
rect 585310 507454 585930 542898
rect 585310 506898 585342 507454
rect 585898 506898 585930 507454
rect 585310 471454 585930 506898
rect 585310 470898 585342 471454
rect 585898 470898 585930 471454
rect 585310 435454 585930 470898
rect 585310 434898 585342 435454
rect 585898 434898 585930 435454
rect 585310 399454 585930 434898
rect 585310 398898 585342 399454
rect 585898 398898 585930 399454
rect 585310 363454 585930 398898
rect 585310 362898 585342 363454
rect 585898 362898 585930 363454
rect 585310 327454 585930 362898
rect 585310 326898 585342 327454
rect 585898 326898 585930 327454
rect 585310 291454 585930 326898
rect 585310 290898 585342 291454
rect 585898 290898 585930 291454
rect 585310 255454 585930 290898
rect 585310 254898 585342 255454
rect 585898 254898 585930 255454
rect 585310 219454 585930 254898
rect 585310 218898 585342 219454
rect 585898 218898 585930 219454
rect 585310 183454 585930 218898
rect 585310 182898 585342 183454
rect 585898 182898 585930 183454
rect 585310 147454 585930 182898
rect 585310 146898 585342 147454
rect 585898 146898 585930 147454
rect 585310 111454 585930 146898
rect 585310 110898 585342 111454
rect 585898 110898 585930 111454
rect 585310 75454 585930 110898
rect 585310 74898 585342 75454
rect 585898 74898 585930 75454
rect 585310 39454 585930 74898
rect 585310 38898 585342 39454
rect 585898 38898 585930 39454
rect 585310 3454 585930 38898
rect 585310 2898 585342 3454
rect 585898 2898 585930 3454
rect 585310 -346 585930 2898
rect 585310 -902 585342 -346
rect 585898 -902 585930 -346
rect 585310 -934 585930 -902
rect 586270 669454 586890 705242
rect 586270 668898 586302 669454
rect 586858 668898 586890 669454
rect 586270 633454 586890 668898
rect 586270 632898 586302 633454
rect 586858 632898 586890 633454
rect 586270 597454 586890 632898
rect 586270 596898 586302 597454
rect 586858 596898 586890 597454
rect 586270 561454 586890 596898
rect 586270 560898 586302 561454
rect 586858 560898 586890 561454
rect 586270 525454 586890 560898
rect 586270 524898 586302 525454
rect 586858 524898 586890 525454
rect 586270 489454 586890 524898
rect 586270 488898 586302 489454
rect 586858 488898 586890 489454
rect 586270 453454 586890 488898
rect 586270 452898 586302 453454
rect 586858 452898 586890 453454
rect 586270 417454 586890 452898
rect 586270 416898 586302 417454
rect 586858 416898 586890 417454
rect 586270 381454 586890 416898
rect 586270 380898 586302 381454
rect 586858 380898 586890 381454
rect 586270 345454 586890 380898
rect 586270 344898 586302 345454
rect 586858 344898 586890 345454
rect 586270 309454 586890 344898
rect 586270 308898 586302 309454
rect 586858 308898 586890 309454
rect 586270 273454 586890 308898
rect 586270 272898 586302 273454
rect 586858 272898 586890 273454
rect 586270 237454 586890 272898
rect 586270 236898 586302 237454
rect 586858 236898 586890 237454
rect 586270 201454 586890 236898
rect 586270 200898 586302 201454
rect 586858 200898 586890 201454
rect 586270 165454 586890 200898
rect 586270 164898 586302 165454
rect 586858 164898 586890 165454
rect 586270 129454 586890 164898
rect 586270 128898 586302 129454
rect 586858 128898 586890 129454
rect 586270 93454 586890 128898
rect 586270 92898 586302 93454
rect 586858 92898 586890 93454
rect 586270 57454 586890 92898
rect 586270 56898 586302 57454
rect 586858 56898 586890 57454
rect 586270 21454 586890 56898
rect 586270 20898 586302 21454
rect 586858 20898 586890 21454
rect 586270 -1306 586890 20898
rect 586270 -1862 586302 -1306
rect 586858 -1862 586890 -1306
rect 586270 -1894 586890 -1862
rect 587230 691174 587850 706202
rect 587230 690618 587262 691174
rect 587818 690618 587850 691174
rect 587230 655174 587850 690618
rect 587230 654618 587262 655174
rect 587818 654618 587850 655174
rect 587230 619174 587850 654618
rect 587230 618618 587262 619174
rect 587818 618618 587850 619174
rect 587230 583174 587850 618618
rect 587230 582618 587262 583174
rect 587818 582618 587850 583174
rect 587230 547174 587850 582618
rect 587230 546618 587262 547174
rect 587818 546618 587850 547174
rect 587230 511174 587850 546618
rect 587230 510618 587262 511174
rect 587818 510618 587850 511174
rect 587230 475174 587850 510618
rect 587230 474618 587262 475174
rect 587818 474618 587850 475174
rect 587230 439174 587850 474618
rect 587230 438618 587262 439174
rect 587818 438618 587850 439174
rect 587230 403174 587850 438618
rect 587230 402618 587262 403174
rect 587818 402618 587850 403174
rect 587230 367174 587850 402618
rect 587230 366618 587262 367174
rect 587818 366618 587850 367174
rect 587230 331174 587850 366618
rect 587230 330618 587262 331174
rect 587818 330618 587850 331174
rect 587230 295174 587850 330618
rect 587230 294618 587262 295174
rect 587818 294618 587850 295174
rect 587230 259174 587850 294618
rect 587230 258618 587262 259174
rect 587818 258618 587850 259174
rect 587230 223174 587850 258618
rect 587230 222618 587262 223174
rect 587818 222618 587850 223174
rect 587230 187174 587850 222618
rect 587230 186618 587262 187174
rect 587818 186618 587850 187174
rect 587230 151174 587850 186618
rect 587230 150618 587262 151174
rect 587818 150618 587850 151174
rect 587230 115174 587850 150618
rect 587230 114618 587262 115174
rect 587818 114618 587850 115174
rect 587230 79174 587850 114618
rect 587230 78618 587262 79174
rect 587818 78618 587850 79174
rect 587230 43174 587850 78618
rect 587230 42618 587262 43174
rect 587818 42618 587850 43174
rect 587230 7174 587850 42618
rect 587230 6618 587262 7174
rect 587818 6618 587850 7174
rect 581514 -2822 581546 -2266
rect 582102 -2822 582134 -2266
rect 581514 -3814 582134 -2822
rect 587230 -2266 587850 6618
rect 587230 -2822 587262 -2266
rect 587818 -2822 587850 -2266
rect 587230 -2854 587850 -2822
rect 588190 673174 588810 707162
rect 588190 672618 588222 673174
rect 588778 672618 588810 673174
rect 588190 637174 588810 672618
rect 588190 636618 588222 637174
rect 588778 636618 588810 637174
rect 588190 601174 588810 636618
rect 588190 600618 588222 601174
rect 588778 600618 588810 601174
rect 588190 565174 588810 600618
rect 588190 564618 588222 565174
rect 588778 564618 588810 565174
rect 588190 529174 588810 564618
rect 588190 528618 588222 529174
rect 588778 528618 588810 529174
rect 588190 493174 588810 528618
rect 588190 492618 588222 493174
rect 588778 492618 588810 493174
rect 588190 457174 588810 492618
rect 588190 456618 588222 457174
rect 588778 456618 588810 457174
rect 588190 421174 588810 456618
rect 588190 420618 588222 421174
rect 588778 420618 588810 421174
rect 588190 385174 588810 420618
rect 588190 384618 588222 385174
rect 588778 384618 588810 385174
rect 588190 349174 588810 384618
rect 588190 348618 588222 349174
rect 588778 348618 588810 349174
rect 588190 313174 588810 348618
rect 588190 312618 588222 313174
rect 588778 312618 588810 313174
rect 588190 277174 588810 312618
rect 588190 276618 588222 277174
rect 588778 276618 588810 277174
rect 588190 241174 588810 276618
rect 588190 240618 588222 241174
rect 588778 240618 588810 241174
rect 588190 205174 588810 240618
rect 588190 204618 588222 205174
rect 588778 204618 588810 205174
rect 588190 169174 588810 204618
rect 588190 168618 588222 169174
rect 588778 168618 588810 169174
rect 588190 133174 588810 168618
rect 588190 132618 588222 133174
rect 588778 132618 588810 133174
rect 588190 97174 588810 132618
rect 588190 96618 588222 97174
rect 588778 96618 588810 97174
rect 588190 61174 588810 96618
rect 588190 60618 588222 61174
rect 588778 60618 588810 61174
rect 588190 25174 588810 60618
rect 588190 24618 588222 25174
rect 588778 24618 588810 25174
rect 588190 -3226 588810 24618
rect 588190 -3782 588222 -3226
rect 588778 -3782 588810 -3226
rect 588190 -3814 588810 -3782
rect 589150 694894 589770 708122
rect 589150 694338 589182 694894
rect 589738 694338 589770 694894
rect 589150 658894 589770 694338
rect 589150 658338 589182 658894
rect 589738 658338 589770 658894
rect 589150 622894 589770 658338
rect 589150 622338 589182 622894
rect 589738 622338 589770 622894
rect 589150 586894 589770 622338
rect 589150 586338 589182 586894
rect 589738 586338 589770 586894
rect 589150 550894 589770 586338
rect 589150 550338 589182 550894
rect 589738 550338 589770 550894
rect 589150 514894 589770 550338
rect 589150 514338 589182 514894
rect 589738 514338 589770 514894
rect 589150 478894 589770 514338
rect 589150 478338 589182 478894
rect 589738 478338 589770 478894
rect 589150 442894 589770 478338
rect 589150 442338 589182 442894
rect 589738 442338 589770 442894
rect 589150 406894 589770 442338
rect 589150 406338 589182 406894
rect 589738 406338 589770 406894
rect 589150 370894 589770 406338
rect 589150 370338 589182 370894
rect 589738 370338 589770 370894
rect 589150 334894 589770 370338
rect 589150 334338 589182 334894
rect 589738 334338 589770 334894
rect 589150 298894 589770 334338
rect 589150 298338 589182 298894
rect 589738 298338 589770 298894
rect 589150 262894 589770 298338
rect 589150 262338 589182 262894
rect 589738 262338 589770 262894
rect 589150 226894 589770 262338
rect 589150 226338 589182 226894
rect 589738 226338 589770 226894
rect 589150 190894 589770 226338
rect 589150 190338 589182 190894
rect 589738 190338 589770 190894
rect 589150 154894 589770 190338
rect 589150 154338 589182 154894
rect 589738 154338 589770 154894
rect 589150 118894 589770 154338
rect 589150 118338 589182 118894
rect 589738 118338 589770 118894
rect 589150 82894 589770 118338
rect 589150 82338 589182 82894
rect 589738 82338 589770 82894
rect 589150 46894 589770 82338
rect 589150 46338 589182 46894
rect 589738 46338 589770 46894
rect 589150 10894 589770 46338
rect 589150 10338 589182 10894
rect 589738 10338 589770 10894
rect 589150 -4186 589770 10338
rect 589150 -4742 589182 -4186
rect 589738 -4742 589770 -4186
rect 589150 -4774 589770 -4742
rect 590110 676894 590730 709082
rect 590110 676338 590142 676894
rect 590698 676338 590730 676894
rect 590110 640894 590730 676338
rect 590110 640338 590142 640894
rect 590698 640338 590730 640894
rect 590110 604894 590730 640338
rect 590110 604338 590142 604894
rect 590698 604338 590730 604894
rect 590110 568894 590730 604338
rect 590110 568338 590142 568894
rect 590698 568338 590730 568894
rect 590110 532894 590730 568338
rect 590110 532338 590142 532894
rect 590698 532338 590730 532894
rect 590110 496894 590730 532338
rect 590110 496338 590142 496894
rect 590698 496338 590730 496894
rect 590110 460894 590730 496338
rect 590110 460338 590142 460894
rect 590698 460338 590730 460894
rect 590110 424894 590730 460338
rect 590110 424338 590142 424894
rect 590698 424338 590730 424894
rect 590110 388894 590730 424338
rect 590110 388338 590142 388894
rect 590698 388338 590730 388894
rect 590110 352894 590730 388338
rect 590110 352338 590142 352894
rect 590698 352338 590730 352894
rect 590110 316894 590730 352338
rect 590110 316338 590142 316894
rect 590698 316338 590730 316894
rect 590110 280894 590730 316338
rect 590110 280338 590142 280894
rect 590698 280338 590730 280894
rect 590110 244894 590730 280338
rect 590110 244338 590142 244894
rect 590698 244338 590730 244894
rect 590110 208894 590730 244338
rect 590110 208338 590142 208894
rect 590698 208338 590730 208894
rect 590110 172894 590730 208338
rect 590110 172338 590142 172894
rect 590698 172338 590730 172894
rect 590110 136894 590730 172338
rect 590110 136338 590142 136894
rect 590698 136338 590730 136894
rect 590110 100894 590730 136338
rect 590110 100338 590142 100894
rect 590698 100338 590730 100894
rect 590110 64894 590730 100338
rect 590110 64338 590142 64894
rect 590698 64338 590730 64894
rect 590110 28894 590730 64338
rect 590110 28338 590142 28894
rect 590698 28338 590730 28894
rect 590110 -5146 590730 28338
rect 590110 -5702 590142 -5146
rect 590698 -5702 590730 -5146
rect 590110 -5734 590730 -5702
rect 591070 698614 591690 710042
rect 591070 698058 591102 698614
rect 591658 698058 591690 698614
rect 591070 662614 591690 698058
rect 591070 662058 591102 662614
rect 591658 662058 591690 662614
rect 591070 626614 591690 662058
rect 591070 626058 591102 626614
rect 591658 626058 591690 626614
rect 591070 590614 591690 626058
rect 591070 590058 591102 590614
rect 591658 590058 591690 590614
rect 591070 554614 591690 590058
rect 591070 554058 591102 554614
rect 591658 554058 591690 554614
rect 591070 518614 591690 554058
rect 591070 518058 591102 518614
rect 591658 518058 591690 518614
rect 591070 482614 591690 518058
rect 591070 482058 591102 482614
rect 591658 482058 591690 482614
rect 591070 446614 591690 482058
rect 591070 446058 591102 446614
rect 591658 446058 591690 446614
rect 591070 410614 591690 446058
rect 591070 410058 591102 410614
rect 591658 410058 591690 410614
rect 591070 374614 591690 410058
rect 591070 374058 591102 374614
rect 591658 374058 591690 374614
rect 591070 338614 591690 374058
rect 591070 338058 591102 338614
rect 591658 338058 591690 338614
rect 591070 302614 591690 338058
rect 591070 302058 591102 302614
rect 591658 302058 591690 302614
rect 591070 266614 591690 302058
rect 591070 266058 591102 266614
rect 591658 266058 591690 266614
rect 591070 230614 591690 266058
rect 591070 230058 591102 230614
rect 591658 230058 591690 230614
rect 591070 194614 591690 230058
rect 591070 194058 591102 194614
rect 591658 194058 591690 194614
rect 591070 158614 591690 194058
rect 591070 158058 591102 158614
rect 591658 158058 591690 158614
rect 591070 122614 591690 158058
rect 591070 122058 591102 122614
rect 591658 122058 591690 122614
rect 591070 86614 591690 122058
rect 591070 86058 591102 86614
rect 591658 86058 591690 86614
rect 591070 50614 591690 86058
rect 591070 50058 591102 50614
rect 591658 50058 591690 50614
rect 591070 14614 591690 50058
rect 591070 14058 591102 14614
rect 591658 14058 591690 14614
rect 591070 -6106 591690 14058
rect 591070 -6662 591102 -6106
rect 591658 -6662 591690 -6106
rect 591070 -6694 591690 -6662
rect 592030 680614 592650 711002
rect 592030 680058 592062 680614
rect 592618 680058 592650 680614
rect 592030 644614 592650 680058
rect 592030 644058 592062 644614
rect 592618 644058 592650 644614
rect 592030 608614 592650 644058
rect 592030 608058 592062 608614
rect 592618 608058 592650 608614
rect 592030 572614 592650 608058
rect 592030 572058 592062 572614
rect 592618 572058 592650 572614
rect 592030 536614 592650 572058
rect 592030 536058 592062 536614
rect 592618 536058 592650 536614
rect 592030 500614 592650 536058
rect 592030 500058 592062 500614
rect 592618 500058 592650 500614
rect 592030 464614 592650 500058
rect 592030 464058 592062 464614
rect 592618 464058 592650 464614
rect 592030 428614 592650 464058
rect 592030 428058 592062 428614
rect 592618 428058 592650 428614
rect 592030 392614 592650 428058
rect 592030 392058 592062 392614
rect 592618 392058 592650 392614
rect 592030 356614 592650 392058
rect 592030 356058 592062 356614
rect 592618 356058 592650 356614
rect 592030 320614 592650 356058
rect 592030 320058 592062 320614
rect 592618 320058 592650 320614
rect 592030 284614 592650 320058
rect 592030 284058 592062 284614
rect 592618 284058 592650 284614
rect 592030 248614 592650 284058
rect 592030 248058 592062 248614
rect 592618 248058 592650 248614
rect 592030 212614 592650 248058
rect 592030 212058 592062 212614
rect 592618 212058 592650 212614
rect 592030 176614 592650 212058
rect 592030 176058 592062 176614
rect 592618 176058 592650 176614
rect 592030 140614 592650 176058
rect 592030 140058 592062 140614
rect 592618 140058 592650 140614
rect 592030 104614 592650 140058
rect 592030 104058 592062 104614
rect 592618 104058 592650 104614
rect 592030 68614 592650 104058
rect 592030 68058 592062 68614
rect 592618 68058 592650 68614
rect 592030 32614 592650 68058
rect 592030 32058 592062 32614
rect 592618 32058 592650 32614
rect 570954 -7622 570986 -7066
rect 571542 -7622 571574 -7066
rect 570954 -7654 571574 -7622
rect 592030 -7066 592650 32058
rect 592030 -7622 592062 -7066
rect 592618 -7622 592650 -7066
rect 592030 -7654 592650 -7622
<< via4 >>
rect -8694 711002 -8138 711558
rect -8694 680058 -8138 680614
rect -8694 644058 -8138 644614
rect -8694 608058 -8138 608614
rect -8694 572058 -8138 572614
rect -8694 536058 -8138 536614
rect -8694 500058 -8138 500614
rect -8694 464058 -8138 464614
rect -8694 428058 -8138 428614
rect -8694 392058 -8138 392614
rect -8694 356058 -8138 356614
rect -8694 320058 -8138 320614
rect -8694 284058 -8138 284614
rect -8694 248058 -8138 248614
rect -8694 212058 -8138 212614
rect -8694 176058 -8138 176614
rect -8694 140058 -8138 140614
rect -8694 104058 -8138 104614
rect -8694 68058 -8138 68614
rect -8694 32058 -8138 32614
rect -7734 710042 -7178 710598
rect 12986 710042 13542 710598
rect -7734 698058 -7178 698614
rect -7734 662058 -7178 662614
rect -7734 626058 -7178 626614
rect -7734 590058 -7178 590614
rect -7734 554058 -7178 554614
rect -7734 518058 -7178 518614
rect -7734 482058 -7178 482614
rect -7734 446058 -7178 446614
rect -7734 410058 -7178 410614
rect -7734 374058 -7178 374614
rect -7734 338058 -7178 338614
rect -7734 302058 -7178 302614
rect -7734 266058 -7178 266614
rect -7734 230058 -7178 230614
rect -7734 194058 -7178 194614
rect -7734 158058 -7178 158614
rect -7734 122058 -7178 122614
rect -7734 86058 -7178 86614
rect -7734 50058 -7178 50614
rect -7734 14058 -7178 14614
rect -6774 709082 -6218 709638
rect -6774 676338 -6218 676894
rect -6774 640338 -6218 640894
rect -6774 604338 -6218 604894
rect -6774 568338 -6218 568894
rect -6774 532338 -6218 532894
rect -6774 496338 -6218 496894
rect -6774 460338 -6218 460894
rect -6774 424338 -6218 424894
rect -6774 388338 -6218 388894
rect -6774 352338 -6218 352894
rect -6774 316338 -6218 316894
rect -6774 280338 -6218 280894
rect -6774 244338 -6218 244894
rect -6774 208338 -6218 208894
rect -6774 172338 -6218 172894
rect -6774 136338 -6218 136894
rect -6774 100338 -6218 100894
rect -6774 64338 -6218 64894
rect -6774 28338 -6218 28894
rect -5814 708122 -5258 708678
rect 9266 708122 9822 708678
rect -5814 694338 -5258 694894
rect -5814 658338 -5258 658894
rect -5814 622338 -5258 622894
rect -5814 586338 -5258 586894
rect -5814 550338 -5258 550894
rect -5814 514338 -5258 514894
rect -5814 478338 -5258 478894
rect -5814 442338 -5258 442894
rect -5814 406338 -5258 406894
rect -5814 370338 -5258 370894
rect -5814 334338 -5258 334894
rect -5814 298338 -5258 298894
rect -5814 262338 -5258 262894
rect -5814 226338 -5258 226894
rect -5814 190338 -5258 190894
rect -5814 154338 -5258 154894
rect -5814 118338 -5258 118894
rect -5814 82338 -5258 82894
rect -5814 46338 -5258 46894
rect -5814 10338 -5258 10894
rect -4854 707162 -4298 707718
rect -4854 672618 -4298 673174
rect -4854 636618 -4298 637174
rect -4854 600618 -4298 601174
rect -4854 564618 -4298 565174
rect -4854 528618 -4298 529174
rect -4854 492618 -4298 493174
rect -4854 456618 -4298 457174
rect -4854 420618 -4298 421174
rect -4854 384618 -4298 385174
rect -4854 348618 -4298 349174
rect -4854 312618 -4298 313174
rect -4854 276618 -4298 277174
rect -4854 240618 -4298 241174
rect -4854 204618 -4298 205174
rect -4854 168618 -4298 169174
rect -4854 132618 -4298 133174
rect -4854 96618 -4298 97174
rect -4854 60618 -4298 61174
rect -4854 24618 -4298 25174
rect -3894 706202 -3338 706758
rect 5546 706202 6102 706758
rect -3894 690618 -3338 691174
rect -3894 654618 -3338 655174
rect -3894 618618 -3338 619174
rect -3894 582618 -3338 583174
rect -3894 546618 -3338 547174
rect -3894 510618 -3338 511174
rect -3894 474618 -3338 475174
rect -3894 438618 -3338 439174
rect -3894 402618 -3338 403174
rect -3894 366618 -3338 367174
rect -3894 330618 -3338 331174
rect -3894 294618 -3338 295174
rect -3894 258618 -3338 259174
rect -3894 222618 -3338 223174
rect -3894 186618 -3338 187174
rect -3894 150618 -3338 151174
rect -3894 114618 -3338 115174
rect -3894 78618 -3338 79174
rect -3894 42618 -3338 43174
rect -3894 6618 -3338 7174
rect -2934 705242 -2378 705798
rect -2934 668898 -2378 669454
rect -2934 632898 -2378 633454
rect -2934 596898 -2378 597454
rect -2934 560898 -2378 561454
rect -2934 524898 -2378 525454
rect -2934 488898 -2378 489454
rect -2934 452898 -2378 453454
rect -2934 416898 -2378 417454
rect -2934 380898 -2378 381454
rect -2934 344898 -2378 345454
rect -2934 308898 -2378 309454
rect -2934 272898 -2378 273454
rect -2934 236898 -2378 237454
rect -2934 200898 -2378 201454
rect -2934 164898 -2378 165454
rect -2934 128898 -2378 129454
rect -2934 92898 -2378 93454
rect -2934 56898 -2378 57454
rect -2934 20898 -2378 21454
rect -1974 704282 -1418 704838
rect -1974 686898 -1418 687454
rect -1974 650898 -1418 651454
rect -1974 614898 -1418 615454
rect -1974 578898 -1418 579454
rect -1974 542898 -1418 543454
rect -1974 506898 -1418 507454
rect -1974 470898 -1418 471454
rect -1974 434898 -1418 435454
rect -1974 398898 -1418 399454
rect -1974 362898 -1418 363454
rect -1974 326898 -1418 327454
rect -1974 290898 -1418 291454
rect -1974 254898 -1418 255454
rect -1974 218898 -1418 219454
rect -1974 182898 -1418 183454
rect -1974 146898 -1418 147454
rect -1974 110898 -1418 111454
rect -1974 74898 -1418 75454
rect -1974 38898 -1418 39454
rect -1974 2898 -1418 3454
rect -1974 -902 -1418 -346
rect 1826 704282 2382 704838
rect 1826 686898 2382 687454
rect 1826 650898 2382 651454
rect 1826 614898 2382 615454
rect 1826 578898 2382 579454
rect 1826 542898 2382 543454
rect 1826 506898 2382 507454
rect 1826 470898 2382 471454
rect 1826 434898 2382 435454
rect 1826 398898 2382 399454
rect 1826 362898 2382 363454
rect 1826 326898 2382 327454
rect 1826 290898 2382 291454
rect 1826 254898 2382 255454
rect 1826 218898 2382 219454
rect 1826 182898 2382 183454
rect 1826 146898 2382 147454
rect 1826 110898 2382 111454
rect 1826 74898 2382 75454
rect 1826 38898 2382 39454
rect 1826 2898 2382 3454
rect 1826 -902 2382 -346
rect -2934 -1862 -2378 -1306
rect 5546 690618 6102 691174
rect 5546 654618 6102 655174
rect 5546 618618 6102 619174
rect 5546 582618 6102 583174
rect 5546 546618 6102 547174
rect 5546 510618 6102 511174
rect 5546 474618 6102 475174
rect 5546 438618 6102 439174
rect 5546 402618 6102 403174
rect 5546 366618 6102 367174
rect 5546 330618 6102 331174
rect 5546 294618 6102 295174
rect 5546 258618 6102 259174
rect 5546 222618 6102 223174
rect 5546 186618 6102 187174
rect 5546 150618 6102 151174
rect 5546 114618 6102 115174
rect 5546 78618 6102 79174
rect 5546 42618 6102 43174
rect 5546 6618 6102 7174
rect -3894 -2822 -3338 -2266
rect 5546 -2822 6102 -2266
rect -4854 -3782 -4298 -3226
rect 9266 694338 9822 694894
rect 9266 658338 9822 658894
rect 9266 622338 9822 622894
rect 9266 586338 9822 586894
rect 9266 550338 9822 550894
rect 9266 514338 9822 514894
rect 9266 478338 9822 478894
rect 9266 442338 9822 442894
rect 9266 406338 9822 406894
rect 9266 370338 9822 370894
rect 9266 334338 9822 334894
rect 9266 298338 9822 298894
rect 9266 262338 9822 262894
rect 9266 226338 9822 226894
rect 9266 190338 9822 190894
rect 9266 154338 9822 154894
rect 9266 118338 9822 118894
rect 9266 82338 9822 82894
rect 9266 46338 9822 46894
rect 9266 10338 9822 10894
rect -5814 -4742 -5258 -4186
rect 9266 -4742 9822 -4186
rect -6774 -5702 -6218 -5146
rect 30986 711002 31542 711558
rect 27266 709082 27822 709638
rect 23546 707162 24102 707718
rect 12986 698058 13542 698614
rect 12986 662058 13542 662614
rect 12986 626058 13542 626614
rect 12986 590058 13542 590614
rect 12986 554058 13542 554614
rect 12986 518058 13542 518614
rect 12986 482058 13542 482614
rect 12986 446058 13542 446614
rect 12986 410058 13542 410614
rect 12986 374058 13542 374614
rect 12986 338058 13542 338614
rect 12986 302058 13542 302614
rect 12986 266058 13542 266614
rect 12986 230058 13542 230614
rect 12986 194058 13542 194614
rect 12986 158058 13542 158614
rect 12986 122058 13542 122614
rect 12986 86058 13542 86614
rect 12986 50058 13542 50614
rect 12986 14058 13542 14614
rect -7734 -6662 -7178 -6106
rect 19826 705242 20382 705798
rect 19826 668898 20382 669454
rect 19826 632898 20382 633454
rect 19826 596898 20382 597454
rect 19826 560898 20382 561454
rect 19826 524898 20382 525454
rect 19826 488898 20382 489454
rect 19826 452898 20382 453454
rect 19826 416898 20382 417454
rect 19826 380898 20382 381454
rect 19826 344898 20382 345454
rect 19826 308898 20382 309454
rect 19826 272898 20382 273454
rect 19826 236898 20382 237454
rect 19826 200898 20382 201454
rect 19826 164898 20382 165454
rect 19826 128898 20382 129454
rect 19826 92898 20382 93454
rect 19826 56898 20382 57454
rect 19826 20898 20382 21454
rect 19826 -1862 20382 -1306
rect 23546 672618 24102 673174
rect 23546 636618 24102 637174
rect 23546 600618 24102 601174
rect 23546 564618 24102 565174
rect 23546 528618 24102 529174
rect 23546 492618 24102 493174
rect 23546 456618 24102 457174
rect 23546 420618 24102 421174
rect 23546 384618 24102 385174
rect 23546 348618 24102 349174
rect 23546 312618 24102 313174
rect 23546 276618 24102 277174
rect 23546 240618 24102 241174
rect 23546 204618 24102 205174
rect 23546 168618 24102 169174
rect 23546 132618 24102 133174
rect 23546 96618 24102 97174
rect 23546 60618 24102 61174
rect 23546 24618 24102 25174
rect 23546 -3782 24102 -3226
rect 27266 676338 27822 676894
rect 27266 640338 27822 640894
rect 27266 604338 27822 604894
rect 27266 568338 27822 568894
rect 27266 532338 27822 532894
rect 27266 496338 27822 496894
rect 27266 460338 27822 460894
rect 27266 424338 27822 424894
rect 27266 388338 27822 388894
rect 27266 352338 27822 352894
rect 27266 316338 27822 316894
rect 27266 280338 27822 280894
rect 27266 244338 27822 244894
rect 27266 208338 27822 208894
rect 27266 172338 27822 172894
rect 27266 136338 27822 136894
rect 27266 100338 27822 100894
rect 27266 64338 27822 64894
rect 27266 28338 27822 28894
rect 27266 -5702 27822 -5146
rect 48986 710042 49542 710598
rect 45266 708122 45822 708678
rect 41546 706202 42102 706758
rect 30986 680058 31542 680614
rect 30986 644058 31542 644614
rect 30986 608058 31542 608614
rect 30986 572058 31542 572614
rect 30986 536058 31542 536614
rect 30986 500058 31542 500614
rect 30986 464058 31542 464614
rect 30986 428058 31542 428614
rect 30986 392058 31542 392614
rect 30986 356058 31542 356614
rect 30986 320058 31542 320614
rect 30986 284058 31542 284614
rect 30986 248058 31542 248614
rect 30986 212058 31542 212614
rect 30986 176058 31542 176614
rect 30986 140058 31542 140614
rect 30986 104058 31542 104614
rect 30986 68058 31542 68614
rect 30986 32058 31542 32614
rect 12986 -6662 13542 -6106
rect -8694 -7622 -8138 -7066
rect 37826 704282 38382 704838
rect 37826 686898 38382 687454
rect 37826 650898 38382 651454
rect 37826 614898 38382 615454
rect 37826 578898 38382 579454
rect 37826 542898 38382 543454
rect 37826 506898 38382 507454
rect 37826 470898 38382 471454
rect 37826 434898 38382 435454
rect 37826 398898 38382 399454
rect 37826 362898 38382 363454
rect 37826 326898 38382 327454
rect 37826 290898 38382 291454
rect 37826 254898 38382 255454
rect 37826 218898 38382 219454
rect 37826 182898 38382 183454
rect 37826 146898 38382 147454
rect 37826 110898 38382 111454
rect 37826 74898 38382 75454
rect 37826 38898 38382 39454
rect 37826 2898 38382 3454
rect 37826 -902 38382 -346
rect 41546 690618 42102 691174
rect 41546 654618 42102 655174
rect 41546 618618 42102 619174
rect 41546 582618 42102 583174
rect 41546 546618 42102 547174
rect 41546 510618 42102 511174
rect 41546 474618 42102 475174
rect 41546 438618 42102 439174
rect 41546 402618 42102 403174
rect 41546 366618 42102 367174
rect 41546 330618 42102 331174
rect 41546 294618 42102 295174
rect 41546 258618 42102 259174
rect 41546 222618 42102 223174
rect 41546 186618 42102 187174
rect 41546 150618 42102 151174
rect 41546 114618 42102 115174
rect 41546 78618 42102 79174
rect 41546 42618 42102 43174
rect 41546 6618 42102 7174
rect 41546 -2822 42102 -2266
rect 45266 694338 45822 694894
rect 45266 658338 45822 658894
rect 45266 622338 45822 622894
rect 45266 586338 45822 586894
rect 45266 550338 45822 550894
rect 45266 514338 45822 514894
rect 45266 478338 45822 478894
rect 45266 442338 45822 442894
rect 45266 406338 45822 406894
rect 45266 370338 45822 370894
rect 45266 334338 45822 334894
rect 45266 298338 45822 298894
rect 45266 262338 45822 262894
rect 45266 226338 45822 226894
rect 45266 190338 45822 190894
rect 45266 154338 45822 154894
rect 45266 118338 45822 118894
rect 45266 82338 45822 82894
rect 45266 46338 45822 46894
rect 45266 10338 45822 10894
rect 45266 -4742 45822 -4186
rect 66986 711002 67542 711558
rect 63266 709082 63822 709638
rect 59546 707162 60102 707718
rect 48986 698058 49542 698614
rect 48986 662058 49542 662614
rect 48986 626058 49542 626614
rect 48986 590058 49542 590614
rect 48986 554058 49542 554614
rect 48986 518058 49542 518614
rect 48986 482058 49542 482614
rect 48986 446058 49542 446614
rect 48986 410058 49542 410614
rect 48986 374058 49542 374614
rect 48986 338058 49542 338614
rect 48986 302058 49542 302614
rect 48986 266058 49542 266614
rect 48986 230058 49542 230614
rect 48986 194058 49542 194614
rect 48986 158058 49542 158614
rect 48986 122058 49542 122614
rect 48986 86058 49542 86614
rect 48986 50058 49542 50614
rect 48986 14058 49542 14614
rect 30986 -7622 31542 -7066
rect 55826 705242 56382 705798
rect 55826 668898 56382 669454
rect 55826 632898 56382 633454
rect 55826 596898 56382 597454
rect 55826 560898 56382 561454
rect 55826 524898 56382 525454
rect 55826 488898 56382 489454
rect 55826 452898 56382 453454
rect 55826 416898 56382 417454
rect 55826 380898 56382 381454
rect 55826 344898 56382 345454
rect 55826 308898 56382 309454
rect 55826 272898 56382 273454
rect 55826 236898 56382 237454
rect 55826 200898 56382 201454
rect 55826 164898 56382 165454
rect 55826 128898 56382 129454
rect 55826 92898 56382 93454
rect 55826 56898 56382 57454
rect 55826 20898 56382 21454
rect 55826 -1862 56382 -1306
rect 59546 672618 60102 673174
rect 59546 636618 60102 637174
rect 59546 600618 60102 601174
rect 59546 564618 60102 565174
rect 59546 528618 60102 529174
rect 59546 492618 60102 493174
rect 59546 456618 60102 457174
rect 59546 420618 60102 421174
rect 59546 384618 60102 385174
rect 59546 348618 60102 349174
rect 59546 312618 60102 313174
rect 59546 276618 60102 277174
rect 59546 240618 60102 241174
rect 59546 204618 60102 205174
rect 59546 168618 60102 169174
rect 59546 132618 60102 133174
rect 59546 96618 60102 97174
rect 59546 60618 60102 61174
rect 59546 24618 60102 25174
rect 59546 -3782 60102 -3226
rect 63266 676338 63822 676894
rect 63266 640338 63822 640894
rect 63266 604338 63822 604894
rect 63266 568338 63822 568894
rect 63266 532338 63822 532894
rect 63266 496338 63822 496894
rect 63266 460338 63822 460894
rect 63266 424338 63822 424894
rect 63266 388338 63822 388894
rect 63266 352338 63822 352894
rect 63266 316338 63822 316894
rect 63266 280338 63822 280894
rect 63266 244338 63822 244894
rect 63266 208338 63822 208894
rect 63266 172338 63822 172894
rect 63266 136338 63822 136894
rect 63266 100338 63822 100894
rect 63266 64338 63822 64894
rect 63266 28338 63822 28894
rect 63266 -5702 63822 -5146
rect 84986 710042 85542 710598
rect 81266 708122 81822 708678
rect 77546 706202 78102 706758
rect 66986 680058 67542 680614
rect 66986 644058 67542 644614
rect 66986 608058 67542 608614
rect 66986 572058 67542 572614
rect 66986 536058 67542 536614
rect 66986 500058 67542 500614
rect 66986 464058 67542 464614
rect 66986 428058 67542 428614
rect 66986 392058 67542 392614
rect 66986 356058 67542 356614
rect 66986 320058 67542 320614
rect 66986 284058 67542 284614
rect 66986 248058 67542 248614
rect 66986 212058 67542 212614
rect 66986 176058 67542 176614
rect 66986 140058 67542 140614
rect 66986 104058 67542 104614
rect 66986 68058 67542 68614
rect 66986 32058 67542 32614
rect 48986 -6662 49542 -6106
rect 73826 704282 74382 704838
rect 73826 686898 74382 687454
rect 73826 650898 74382 651454
rect 73826 614898 74382 615454
rect 73826 578898 74382 579454
rect 73826 542898 74382 543454
rect 73826 506898 74382 507454
rect 73826 470898 74382 471454
rect 73826 434898 74382 435454
rect 73826 398898 74382 399454
rect 73826 362898 74382 363454
rect 73826 326898 74382 327454
rect 73826 290898 74382 291454
rect 73826 254898 74382 255454
rect 73826 218898 74382 219454
rect 73826 182898 74382 183454
rect 73826 146898 74382 147454
rect 73826 110898 74382 111454
rect 73826 74898 74382 75454
rect 73826 38898 74382 39454
rect 73826 2898 74382 3454
rect 73826 -902 74382 -346
rect 77546 690618 78102 691174
rect 77546 654618 78102 655174
rect 77546 618618 78102 619174
rect 77546 582618 78102 583174
rect 77546 546618 78102 547174
rect 77546 510618 78102 511174
rect 77546 474618 78102 475174
rect 77546 438618 78102 439174
rect 77546 402618 78102 403174
rect 77546 366618 78102 367174
rect 77546 330618 78102 331174
rect 77546 294618 78102 295174
rect 77546 258618 78102 259174
rect 77546 222618 78102 223174
rect 77546 186618 78102 187174
rect 77546 150618 78102 151174
rect 77546 114618 78102 115174
rect 77546 78618 78102 79174
rect 77546 42618 78102 43174
rect 77546 6618 78102 7174
rect 77546 -2822 78102 -2266
rect 81266 694338 81822 694894
rect 81266 658338 81822 658894
rect 81266 622338 81822 622894
rect 81266 586338 81822 586894
rect 81266 550338 81822 550894
rect 81266 514338 81822 514894
rect 81266 478338 81822 478894
rect 81266 442338 81822 442894
rect 81266 406338 81822 406894
rect 81266 370338 81822 370894
rect 81266 334338 81822 334894
rect 81266 298338 81822 298894
rect 81266 262338 81822 262894
rect 81266 226338 81822 226894
rect 81266 190338 81822 190894
rect 81266 154338 81822 154894
rect 81266 118338 81822 118894
rect 81266 82338 81822 82894
rect 81266 46338 81822 46894
rect 81266 10338 81822 10894
rect 81266 -4742 81822 -4186
rect 102986 711002 103542 711558
rect 99266 709082 99822 709638
rect 95546 707162 96102 707718
rect 84986 698058 85542 698614
rect 84986 662058 85542 662614
rect 84986 626058 85542 626614
rect 84986 590058 85542 590614
rect 84986 554058 85542 554614
rect 84986 518058 85542 518614
rect 84986 482058 85542 482614
rect 84986 446058 85542 446614
rect 84986 410058 85542 410614
rect 84986 374058 85542 374614
rect 84986 338058 85542 338614
rect 84986 302058 85542 302614
rect 84986 266058 85542 266614
rect 84986 230058 85542 230614
rect 84986 194058 85542 194614
rect 84986 158058 85542 158614
rect 84986 122058 85542 122614
rect 84986 86058 85542 86614
rect 84986 50058 85542 50614
rect 84986 14058 85542 14614
rect 66986 -7622 67542 -7066
rect 91826 705242 92382 705798
rect 91826 668898 92382 669454
rect 91826 632898 92382 633454
rect 91826 596898 92382 597454
rect 91826 560898 92382 561454
rect 91826 524898 92382 525454
rect 91826 488898 92382 489454
rect 91826 452898 92382 453454
rect 91826 416898 92382 417454
rect 91826 380898 92382 381454
rect 91826 344898 92382 345454
rect 91826 308898 92382 309454
rect 91826 272898 92382 273454
rect 91826 236898 92382 237454
rect 91826 200898 92382 201454
rect 91826 164898 92382 165454
rect 91826 128898 92382 129454
rect 91826 92898 92382 93454
rect 91826 56898 92382 57454
rect 91826 20898 92382 21454
rect 91826 -1862 92382 -1306
rect 95546 672618 96102 673174
rect 95546 636618 96102 637174
rect 95546 600618 96102 601174
rect 95546 564618 96102 565174
rect 95546 528618 96102 529174
rect 95546 492618 96102 493174
rect 95546 456618 96102 457174
rect 95546 420618 96102 421174
rect 95546 384618 96102 385174
rect 95546 348618 96102 349174
rect 95546 312618 96102 313174
rect 95546 276618 96102 277174
rect 95546 240618 96102 241174
rect 95546 204618 96102 205174
rect 95546 168618 96102 169174
rect 95546 132618 96102 133174
rect 95546 96618 96102 97174
rect 95546 60618 96102 61174
rect 95546 24618 96102 25174
rect 95546 -3782 96102 -3226
rect 99266 676338 99822 676894
rect 99266 640338 99822 640894
rect 99266 604338 99822 604894
rect 99266 568338 99822 568894
rect 99266 532338 99822 532894
rect 99266 496338 99822 496894
rect 99266 460338 99822 460894
rect 99266 424338 99822 424894
rect 99266 388338 99822 388894
rect 99266 352338 99822 352894
rect 99266 316338 99822 316894
rect 99266 280338 99822 280894
rect 99266 244338 99822 244894
rect 99266 208338 99822 208894
rect 99266 172338 99822 172894
rect 99266 136338 99822 136894
rect 99266 100338 99822 100894
rect 99266 64338 99822 64894
rect 99266 28338 99822 28894
rect 99266 -5702 99822 -5146
rect 120986 710042 121542 710598
rect 117266 708122 117822 708678
rect 113546 706202 114102 706758
rect 102986 680058 103542 680614
rect 102986 644058 103542 644614
rect 102986 608058 103542 608614
rect 102986 572058 103542 572614
rect 102986 536058 103542 536614
rect 102986 500058 103542 500614
rect 102986 464058 103542 464614
rect 102986 428058 103542 428614
rect 102986 392058 103542 392614
rect 102986 356058 103542 356614
rect 102986 320058 103542 320614
rect 102986 284058 103542 284614
rect 102986 248058 103542 248614
rect 102986 212058 103542 212614
rect 102986 176058 103542 176614
rect 102986 140058 103542 140614
rect 102986 104058 103542 104614
rect 102986 68058 103542 68614
rect 102986 32058 103542 32614
rect 84986 -6662 85542 -6106
rect 109826 704282 110382 704838
rect 109826 686898 110382 687454
rect 109826 650898 110382 651454
rect 109826 614898 110382 615454
rect 109826 578898 110382 579454
rect 109826 542898 110382 543454
rect 109826 506898 110382 507454
rect 109826 470898 110382 471454
rect 109826 434898 110382 435454
rect 109826 398898 110382 399454
rect 109826 362898 110382 363454
rect 109826 326898 110382 327454
rect 109826 290898 110382 291454
rect 109826 254898 110382 255454
rect 109826 218898 110382 219454
rect 109826 182898 110382 183454
rect 109826 146898 110382 147454
rect 109826 110898 110382 111454
rect 109826 74898 110382 75454
rect 109826 38898 110382 39454
rect 109826 2898 110382 3454
rect 109826 -902 110382 -346
rect 113546 690618 114102 691174
rect 113546 654618 114102 655174
rect 113546 618618 114102 619174
rect 113546 582618 114102 583174
rect 113546 546618 114102 547174
rect 113546 510618 114102 511174
rect 113546 474618 114102 475174
rect 113546 438618 114102 439174
rect 113546 402618 114102 403174
rect 113546 366618 114102 367174
rect 113546 330618 114102 331174
rect 113546 294618 114102 295174
rect 113546 258618 114102 259174
rect 113546 222618 114102 223174
rect 113546 186618 114102 187174
rect 113546 150618 114102 151174
rect 113546 114618 114102 115174
rect 113546 78618 114102 79174
rect 113546 42618 114102 43174
rect 113546 6618 114102 7174
rect 113546 -2822 114102 -2266
rect 117266 694338 117822 694894
rect 117266 658338 117822 658894
rect 117266 622338 117822 622894
rect 117266 586338 117822 586894
rect 117266 550338 117822 550894
rect 117266 514338 117822 514894
rect 117266 478338 117822 478894
rect 117266 442338 117822 442894
rect 117266 406338 117822 406894
rect 117266 370338 117822 370894
rect 117266 334338 117822 334894
rect 117266 298338 117822 298894
rect 117266 262338 117822 262894
rect 117266 226338 117822 226894
rect 117266 190338 117822 190894
rect 117266 154338 117822 154894
rect 117266 118338 117822 118894
rect 117266 82338 117822 82894
rect 117266 46338 117822 46894
rect 117266 10338 117822 10894
rect 117266 -4742 117822 -4186
rect 138986 711002 139542 711558
rect 135266 709082 135822 709638
rect 131546 707162 132102 707718
rect 120986 698058 121542 698614
rect 120986 662058 121542 662614
rect 120986 626058 121542 626614
rect 120986 590058 121542 590614
rect 120986 554058 121542 554614
rect 120986 518058 121542 518614
rect 120986 482058 121542 482614
rect 120986 446058 121542 446614
rect 120986 410058 121542 410614
rect 120986 374058 121542 374614
rect 120986 338058 121542 338614
rect 120986 302058 121542 302614
rect 120986 266058 121542 266614
rect 120986 230058 121542 230614
rect 120986 194058 121542 194614
rect 120986 158058 121542 158614
rect 120986 122058 121542 122614
rect 120986 86058 121542 86614
rect 120986 50058 121542 50614
rect 120986 14058 121542 14614
rect 102986 -7622 103542 -7066
rect 127826 705242 128382 705798
rect 127826 668898 128382 669454
rect 127826 632898 128382 633454
rect 127826 596898 128382 597454
rect 127826 560898 128382 561454
rect 127826 524898 128382 525454
rect 127826 488898 128382 489454
rect 127826 452898 128382 453454
rect 127826 416898 128382 417454
rect 127826 380898 128382 381454
rect 127826 344898 128382 345454
rect 127826 308898 128382 309454
rect 127826 272898 128382 273454
rect 127826 236898 128382 237454
rect 127826 200898 128382 201454
rect 127826 164898 128382 165454
rect 127826 128898 128382 129454
rect 127826 92898 128382 93454
rect 127826 56898 128382 57454
rect 127826 20898 128382 21454
rect 127826 -1862 128382 -1306
rect 131546 672618 132102 673174
rect 131546 636618 132102 637174
rect 131546 600618 132102 601174
rect 131546 564618 132102 565174
rect 131546 528618 132102 529174
rect 131546 492618 132102 493174
rect 131546 456618 132102 457174
rect 131546 420618 132102 421174
rect 131546 384618 132102 385174
rect 131546 348618 132102 349174
rect 131546 312618 132102 313174
rect 131546 276618 132102 277174
rect 131546 240618 132102 241174
rect 131546 204618 132102 205174
rect 131546 168618 132102 169174
rect 131546 132618 132102 133174
rect 131546 96618 132102 97174
rect 131546 60618 132102 61174
rect 131546 24618 132102 25174
rect 131546 -3782 132102 -3226
rect 135266 676338 135822 676894
rect 135266 640338 135822 640894
rect 135266 604338 135822 604894
rect 135266 568338 135822 568894
rect 135266 532338 135822 532894
rect 135266 496338 135822 496894
rect 135266 460338 135822 460894
rect 135266 424338 135822 424894
rect 135266 388338 135822 388894
rect 135266 352338 135822 352894
rect 135266 316338 135822 316894
rect 135266 280338 135822 280894
rect 135266 244338 135822 244894
rect 135266 208338 135822 208894
rect 135266 172338 135822 172894
rect 135266 136338 135822 136894
rect 135266 100338 135822 100894
rect 135266 64338 135822 64894
rect 135266 28338 135822 28894
rect 135266 -5702 135822 -5146
rect 156986 710042 157542 710598
rect 153266 708122 153822 708678
rect 149546 706202 150102 706758
rect 138986 680058 139542 680614
rect 138986 644058 139542 644614
rect 138986 608058 139542 608614
rect 138986 572058 139542 572614
rect 138986 536058 139542 536614
rect 138986 500058 139542 500614
rect 138986 464058 139542 464614
rect 138986 428058 139542 428614
rect 138986 392058 139542 392614
rect 138986 356058 139542 356614
rect 138986 320058 139542 320614
rect 138986 284058 139542 284614
rect 138986 248058 139542 248614
rect 138986 212058 139542 212614
rect 138986 176058 139542 176614
rect 138986 140058 139542 140614
rect 138986 104058 139542 104614
rect 138986 68058 139542 68614
rect 138986 32058 139542 32614
rect 120986 -6662 121542 -6106
rect 145826 704282 146382 704838
rect 145826 686898 146382 687454
rect 145826 650898 146382 651454
rect 145826 614898 146382 615454
rect 145826 578898 146382 579454
rect 145826 542898 146382 543454
rect 145826 506898 146382 507454
rect 145826 470898 146382 471454
rect 145826 434898 146382 435454
rect 145826 398898 146382 399454
rect 145826 362898 146382 363454
rect 145826 326898 146382 327454
rect 145826 290898 146382 291454
rect 145826 254898 146382 255454
rect 145826 218898 146382 219454
rect 145826 182898 146382 183454
rect 145826 146898 146382 147454
rect 145826 110898 146382 111454
rect 145826 74898 146382 75454
rect 145826 38898 146382 39454
rect 145826 2898 146382 3454
rect 145826 -902 146382 -346
rect 149546 690618 150102 691174
rect 149546 654618 150102 655174
rect 149546 618618 150102 619174
rect 149546 582618 150102 583174
rect 149546 546618 150102 547174
rect 149546 510618 150102 511174
rect 149546 474618 150102 475174
rect 149546 438618 150102 439174
rect 149546 402618 150102 403174
rect 149546 366618 150102 367174
rect 149546 330618 150102 331174
rect 149546 294618 150102 295174
rect 149546 258618 150102 259174
rect 149546 222618 150102 223174
rect 149546 186618 150102 187174
rect 149546 150618 150102 151174
rect 149546 114618 150102 115174
rect 149546 78618 150102 79174
rect 149546 42618 150102 43174
rect 149546 6618 150102 7174
rect 149546 -2822 150102 -2266
rect 153266 694338 153822 694894
rect 153266 658338 153822 658894
rect 153266 622338 153822 622894
rect 153266 586338 153822 586894
rect 153266 550338 153822 550894
rect 153266 514338 153822 514894
rect 153266 478338 153822 478894
rect 153266 442338 153822 442894
rect 153266 406338 153822 406894
rect 153266 370338 153822 370894
rect 153266 334338 153822 334894
rect 153266 298338 153822 298894
rect 153266 262338 153822 262894
rect 153266 226338 153822 226894
rect 153266 190338 153822 190894
rect 153266 154338 153822 154894
rect 153266 118338 153822 118894
rect 153266 82338 153822 82894
rect 153266 46338 153822 46894
rect 153266 10338 153822 10894
rect 153266 -4742 153822 -4186
rect 174986 711002 175542 711558
rect 171266 709082 171822 709638
rect 167546 707162 168102 707718
rect 156986 698058 157542 698614
rect 156986 662058 157542 662614
rect 156986 626058 157542 626614
rect 156986 590058 157542 590614
rect 156986 554058 157542 554614
rect 156986 518058 157542 518614
rect 156986 482058 157542 482614
rect 156986 446058 157542 446614
rect 156986 410058 157542 410614
rect 156986 374058 157542 374614
rect 156986 338058 157542 338614
rect 156986 302058 157542 302614
rect 156986 266058 157542 266614
rect 156986 230058 157542 230614
rect 156986 194058 157542 194614
rect 156986 158058 157542 158614
rect 156986 122058 157542 122614
rect 156986 86058 157542 86614
rect 156986 50058 157542 50614
rect 156986 14058 157542 14614
rect 138986 -7622 139542 -7066
rect 163826 705242 164382 705798
rect 163826 668898 164382 669454
rect 163826 632898 164382 633454
rect 163826 596898 164382 597454
rect 163826 560898 164382 561454
rect 163826 524898 164382 525454
rect 163826 488898 164382 489454
rect 163826 452898 164382 453454
rect 163826 416898 164382 417454
rect 163826 380898 164382 381454
rect 163826 344898 164382 345454
rect 163826 308898 164382 309454
rect 163826 272898 164382 273454
rect 163826 236898 164382 237454
rect 163826 200898 164382 201454
rect 163826 164898 164382 165454
rect 163826 128898 164382 129454
rect 163826 92898 164382 93454
rect 163826 56898 164382 57454
rect 163826 20898 164382 21454
rect 163826 -1862 164382 -1306
rect 167546 672618 168102 673174
rect 167546 636618 168102 637174
rect 167546 600618 168102 601174
rect 167546 564618 168102 565174
rect 167546 528618 168102 529174
rect 167546 492618 168102 493174
rect 167546 456618 168102 457174
rect 167546 420618 168102 421174
rect 167546 384618 168102 385174
rect 167546 348618 168102 349174
rect 167546 312618 168102 313174
rect 167546 276618 168102 277174
rect 167546 240618 168102 241174
rect 167546 204618 168102 205174
rect 167546 168618 168102 169174
rect 167546 132618 168102 133174
rect 167546 96618 168102 97174
rect 167546 60618 168102 61174
rect 167546 24618 168102 25174
rect 167546 -3782 168102 -3226
rect 171266 676338 171822 676894
rect 171266 640338 171822 640894
rect 171266 604338 171822 604894
rect 171266 568338 171822 568894
rect 171266 532338 171822 532894
rect 171266 496338 171822 496894
rect 171266 460338 171822 460894
rect 171266 424338 171822 424894
rect 171266 388338 171822 388894
rect 171266 352338 171822 352894
rect 171266 316338 171822 316894
rect 171266 280338 171822 280894
rect 171266 244338 171822 244894
rect 171266 208338 171822 208894
rect 171266 172338 171822 172894
rect 171266 136338 171822 136894
rect 171266 100338 171822 100894
rect 171266 64338 171822 64894
rect 171266 28338 171822 28894
rect 171266 -5702 171822 -5146
rect 192986 710042 193542 710598
rect 189266 708122 189822 708678
rect 185546 706202 186102 706758
rect 174986 680058 175542 680614
rect 174986 644058 175542 644614
rect 174986 608058 175542 608614
rect 174986 572058 175542 572614
rect 174986 536058 175542 536614
rect 174986 500058 175542 500614
rect 174986 464058 175542 464614
rect 174986 428058 175542 428614
rect 174986 392058 175542 392614
rect 174986 356058 175542 356614
rect 174986 320058 175542 320614
rect 174986 284058 175542 284614
rect 174986 248058 175542 248614
rect 174986 212058 175542 212614
rect 174986 176058 175542 176614
rect 174986 140058 175542 140614
rect 174986 104058 175542 104614
rect 174986 68058 175542 68614
rect 174986 32058 175542 32614
rect 156986 -6662 157542 -6106
rect 181826 704282 182382 704838
rect 181826 686898 182382 687454
rect 181826 650898 182382 651454
rect 181826 614898 182382 615454
rect 181826 578898 182382 579454
rect 181826 542898 182382 543454
rect 181826 506898 182382 507454
rect 181826 470898 182382 471454
rect 181826 434898 182382 435454
rect 181826 398898 182382 399454
rect 181826 362898 182382 363454
rect 181826 326898 182382 327454
rect 181826 290898 182382 291454
rect 181826 254898 182382 255454
rect 181826 218898 182382 219454
rect 181826 182898 182382 183454
rect 181826 146898 182382 147454
rect 181826 110898 182382 111454
rect 181826 74898 182382 75454
rect 181826 38898 182382 39454
rect 181826 2898 182382 3454
rect 181826 -902 182382 -346
rect 185546 690618 186102 691174
rect 185546 654618 186102 655174
rect 185546 618618 186102 619174
rect 185546 582618 186102 583174
rect 185546 546618 186102 547174
rect 185546 510618 186102 511174
rect 185546 474618 186102 475174
rect 185546 438618 186102 439174
rect 185546 402618 186102 403174
rect 185546 366618 186102 367174
rect 185546 330618 186102 331174
rect 185546 294618 186102 295174
rect 185546 258618 186102 259174
rect 185546 222618 186102 223174
rect 185546 186618 186102 187174
rect 185546 150618 186102 151174
rect 185546 114618 186102 115174
rect 185546 78618 186102 79174
rect 185546 42618 186102 43174
rect 185546 6618 186102 7174
rect 185546 -2822 186102 -2266
rect 189266 694338 189822 694894
rect 189266 658338 189822 658894
rect 189266 622338 189822 622894
rect 189266 586338 189822 586894
rect 189266 550338 189822 550894
rect 189266 514338 189822 514894
rect 189266 478338 189822 478894
rect 189266 442338 189822 442894
rect 189266 406338 189822 406894
rect 189266 370338 189822 370894
rect 189266 334338 189822 334894
rect 189266 298338 189822 298894
rect 189266 262338 189822 262894
rect 189266 226338 189822 226894
rect 189266 190338 189822 190894
rect 189266 154338 189822 154894
rect 189266 118338 189822 118894
rect 189266 82338 189822 82894
rect 189266 46338 189822 46894
rect 189266 10338 189822 10894
rect 189266 -4742 189822 -4186
rect 210986 711002 211542 711558
rect 207266 709082 207822 709638
rect 203546 707162 204102 707718
rect 192986 698058 193542 698614
rect 192986 662058 193542 662614
rect 192986 626058 193542 626614
rect 192986 590058 193542 590614
rect 192986 554058 193542 554614
rect 192986 518058 193542 518614
rect 192986 482058 193542 482614
rect 192986 446058 193542 446614
rect 192986 410058 193542 410614
rect 192986 374058 193542 374614
rect 192986 338058 193542 338614
rect 192986 302058 193542 302614
rect 192986 266058 193542 266614
rect 192986 230058 193542 230614
rect 192986 194058 193542 194614
rect 192986 158058 193542 158614
rect 192986 122058 193542 122614
rect 192986 86058 193542 86614
rect 192986 50058 193542 50614
rect 192986 14058 193542 14614
rect 174986 -7622 175542 -7066
rect 199826 705242 200382 705798
rect 199826 668898 200382 669454
rect 199826 632898 200382 633454
rect 199826 596898 200382 597454
rect 199826 560898 200382 561454
rect 199826 524898 200382 525454
rect 199826 488898 200382 489454
rect 199826 452898 200382 453454
rect 199826 416898 200382 417454
rect 199826 380898 200382 381454
rect 199826 344898 200382 345454
rect 199826 308898 200382 309454
rect 199826 272898 200382 273454
rect 199826 236898 200382 237454
rect 199826 200898 200382 201454
rect 199826 164898 200382 165454
rect 199826 128898 200382 129454
rect 199826 92898 200382 93454
rect 199826 56898 200382 57454
rect 199826 20898 200382 21454
rect 199826 -1862 200382 -1306
rect 203546 672618 204102 673174
rect 203546 636618 204102 637174
rect 203546 600618 204102 601174
rect 203546 564618 204102 565174
rect 203546 528618 204102 529174
rect 203546 492618 204102 493174
rect 203546 456618 204102 457174
rect 203546 420618 204102 421174
rect 203546 384618 204102 385174
rect 203546 348618 204102 349174
rect 203546 312618 204102 313174
rect 203546 276618 204102 277174
rect 203546 240618 204102 241174
rect 203546 204618 204102 205174
rect 203546 168618 204102 169174
rect 203546 132618 204102 133174
rect 203546 96618 204102 97174
rect 203546 60618 204102 61174
rect 203546 24618 204102 25174
rect 203546 -3782 204102 -3226
rect 207266 676338 207822 676894
rect 207266 640338 207822 640894
rect 207266 604338 207822 604894
rect 207266 568338 207822 568894
rect 207266 532338 207822 532894
rect 207266 496338 207822 496894
rect 207266 460338 207822 460894
rect 207266 424338 207822 424894
rect 207266 388338 207822 388894
rect 207266 352338 207822 352894
rect 207266 316338 207822 316894
rect 207266 280338 207822 280894
rect 207266 244338 207822 244894
rect 207266 208338 207822 208894
rect 207266 172338 207822 172894
rect 207266 136338 207822 136894
rect 207266 100338 207822 100894
rect 207266 64338 207822 64894
rect 207266 28338 207822 28894
rect 207266 -5702 207822 -5146
rect 228986 710042 229542 710598
rect 225266 708122 225822 708678
rect 221546 706202 222102 706758
rect 210986 680058 211542 680614
rect 210986 644058 211542 644614
rect 210986 608058 211542 608614
rect 210986 572058 211542 572614
rect 210986 536058 211542 536614
rect 210986 500058 211542 500614
rect 210986 464058 211542 464614
rect 210986 428058 211542 428614
rect 210986 392058 211542 392614
rect 210986 356058 211542 356614
rect 210986 320058 211542 320614
rect 210986 284058 211542 284614
rect 210986 248058 211542 248614
rect 210986 212058 211542 212614
rect 210986 176058 211542 176614
rect 210986 140058 211542 140614
rect 210986 104058 211542 104614
rect 210986 68058 211542 68614
rect 210986 32058 211542 32614
rect 192986 -6662 193542 -6106
rect 217826 704282 218382 704838
rect 217826 686898 218382 687454
rect 217826 650898 218382 651454
rect 217826 614898 218382 615454
rect 217826 578898 218382 579454
rect 217826 542898 218382 543454
rect 217826 506898 218382 507454
rect 217826 470898 218382 471454
rect 217826 434898 218382 435454
rect 217826 398898 218382 399454
rect 217826 362898 218382 363454
rect 217826 326898 218382 327454
rect 217826 290898 218382 291454
rect 217826 254898 218382 255454
rect 217826 218898 218382 219454
rect 217826 182898 218382 183454
rect 217826 146898 218382 147454
rect 217826 110898 218382 111454
rect 217826 74898 218382 75454
rect 217826 38898 218382 39454
rect 217826 2898 218382 3454
rect 217826 -902 218382 -346
rect 221546 690618 222102 691174
rect 221546 654618 222102 655174
rect 221546 618618 222102 619174
rect 221546 582618 222102 583174
rect 221546 546618 222102 547174
rect 221546 510618 222102 511174
rect 221546 474618 222102 475174
rect 221546 438618 222102 439174
rect 221546 402618 222102 403174
rect 221546 366618 222102 367174
rect 221546 330618 222102 331174
rect 221546 294618 222102 295174
rect 221546 258618 222102 259174
rect 221546 222618 222102 223174
rect 221546 186618 222102 187174
rect 221546 150618 222102 151174
rect 221546 114618 222102 115174
rect 221546 78618 222102 79174
rect 221546 42618 222102 43174
rect 221546 6618 222102 7174
rect 221546 -2822 222102 -2266
rect 225266 694338 225822 694894
rect 225266 658338 225822 658894
rect 225266 622338 225822 622894
rect 225266 586338 225822 586894
rect 225266 550338 225822 550894
rect 225266 514338 225822 514894
rect 225266 478338 225822 478894
rect 225266 442338 225822 442894
rect 225266 406338 225822 406894
rect 225266 370338 225822 370894
rect 225266 334338 225822 334894
rect 225266 298338 225822 298894
rect 225266 262338 225822 262894
rect 225266 226338 225822 226894
rect 225266 190338 225822 190894
rect 225266 154338 225822 154894
rect 225266 118338 225822 118894
rect 225266 82338 225822 82894
rect 225266 46338 225822 46894
rect 225266 10338 225822 10894
rect 225266 -4742 225822 -4186
rect 246986 711002 247542 711558
rect 243266 709082 243822 709638
rect 239546 707162 240102 707718
rect 228986 698058 229542 698614
rect 228986 662058 229542 662614
rect 228986 626058 229542 626614
rect 228986 590058 229542 590614
rect 228986 554058 229542 554614
rect 228986 518058 229542 518614
rect 235826 705242 236382 705798
rect 235826 668898 236382 669454
rect 235826 632898 236382 633454
rect 235826 596898 236382 597454
rect 235826 560898 236382 561454
rect 235826 524898 236382 525454
rect 239546 672618 240102 673174
rect 239546 636618 240102 637174
rect 239546 600618 240102 601174
rect 239546 564618 240102 565174
rect 239546 528618 240102 529174
rect 239546 492618 240102 493174
rect 243266 676338 243822 676894
rect 243266 640338 243822 640894
rect 243266 604338 243822 604894
rect 243266 568338 243822 568894
rect 243266 532338 243822 532894
rect 243266 496338 243822 496894
rect 264986 710042 265542 710598
rect 261266 708122 261822 708678
rect 257546 706202 258102 706758
rect 246986 680058 247542 680614
rect 246986 644058 247542 644614
rect 246986 608058 247542 608614
rect 246986 572058 247542 572614
rect 246986 536058 247542 536614
rect 246986 500058 247542 500614
rect 253826 704282 254382 704838
rect 253826 686898 254382 687454
rect 253826 650898 254382 651454
rect 253826 614898 254382 615454
rect 253826 578898 254382 579454
rect 253826 542898 254382 543454
rect 253826 506898 254382 507454
rect 257546 690618 258102 691174
rect 257546 654618 258102 655174
rect 257546 618618 258102 619174
rect 257546 582618 258102 583174
rect 257546 546618 258102 547174
rect 257546 510618 258102 511174
rect 261266 694338 261822 694894
rect 261266 658338 261822 658894
rect 261266 622338 261822 622894
rect 261266 586338 261822 586894
rect 261266 550338 261822 550894
rect 261266 514338 261822 514894
rect 282986 711002 283542 711558
rect 279266 709082 279822 709638
rect 275546 707162 276102 707718
rect 264986 698058 265542 698614
rect 264986 662058 265542 662614
rect 264986 626058 265542 626614
rect 264986 590058 265542 590614
rect 264986 554058 265542 554614
rect 264986 518058 265542 518614
rect 271826 705242 272382 705798
rect 271826 668898 272382 669454
rect 271826 632898 272382 633454
rect 271826 596898 272382 597454
rect 271826 560898 272382 561454
rect 271826 524898 272382 525454
rect 275546 672618 276102 673174
rect 275546 636618 276102 637174
rect 275546 600618 276102 601174
rect 275546 564618 276102 565174
rect 275546 528618 276102 529174
rect 275546 492618 276102 493174
rect 279266 676338 279822 676894
rect 279266 640338 279822 640894
rect 279266 604338 279822 604894
rect 279266 568338 279822 568894
rect 279266 532338 279822 532894
rect 279266 496338 279822 496894
rect 300986 710042 301542 710598
rect 297266 708122 297822 708678
rect 293546 706202 294102 706758
rect 282986 680058 283542 680614
rect 282986 644058 283542 644614
rect 282986 608058 283542 608614
rect 282986 572058 283542 572614
rect 282986 536058 283542 536614
rect 282986 500058 283542 500614
rect 289826 704282 290382 704838
rect 289826 686898 290382 687454
rect 289826 650898 290382 651454
rect 289826 614898 290382 615454
rect 289826 578898 290382 579454
rect 289826 542898 290382 543454
rect 289826 506898 290382 507454
rect 293546 690618 294102 691174
rect 293546 654618 294102 655174
rect 293546 618618 294102 619174
rect 293546 582618 294102 583174
rect 293546 546618 294102 547174
rect 293546 510618 294102 511174
rect 297266 694338 297822 694894
rect 297266 658338 297822 658894
rect 297266 622338 297822 622894
rect 297266 586338 297822 586894
rect 297266 550338 297822 550894
rect 297266 514338 297822 514894
rect 318986 711002 319542 711558
rect 315266 709082 315822 709638
rect 311546 707162 312102 707718
rect 300986 698058 301542 698614
rect 300986 662058 301542 662614
rect 300986 626058 301542 626614
rect 300986 590058 301542 590614
rect 300986 554058 301542 554614
rect 300986 518058 301542 518614
rect 307826 705242 308382 705798
rect 307826 668898 308382 669454
rect 307826 632898 308382 633454
rect 307826 596898 308382 597454
rect 307826 560898 308382 561454
rect 307826 524898 308382 525454
rect 311546 672618 312102 673174
rect 311546 636618 312102 637174
rect 311546 600618 312102 601174
rect 311546 564618 312102 565174
rect 311546 528618 312102 529174
rect 311546 492618 312102 493174
rect 315266 676338 315822 676894
rect 315266 640338 315822 640894
rect 315266 604338 315822 604894
rect 315266 568338 315822 568894
rect 315266 532338 315822 532894
rect 315266 496338 315822 496894
rect 336986 710042 337542 710598
rect 333266 708122 333822 708678
rect 329546 706202 330102 706758
rect 318986 680058 319542 680614
rect 318986 644058 319542 644614
rect 318986 608058 319542 608614
rect 318986 572058 319542 572614
rect 318986 536058 319542 536614
rect 318986 500058 319542 500614
rect 325826 704282 326382 704838
rect 325826 686898 326382 687454
rect 325826 650898 326382 651454
rect 325826 614898 326382 615454
rect 325826 578898 326382 579454
rect 325826 542898 326382 543454
rect 325826 506898 326382 507454
rect 329546 690618 330102 691174
rect 329546 654618 330102 655174
rect 329546 618618 330102 619174
rect 329546 582618 330102 583174
rect 329546 546618 330102 547174
rect 329546 510618 330102 511174
rect 333266 694338 333822 694894
rect 333266 658338 333822 658894
rect 333266 622338 333822 622894
rect 333266 586338 333822 586894
rect 333266 550338 333822 550894
rect 333266 514338 333822 514894
rect 354986 711002 355542 711558
rect 351266 709082 351822 709638
rect 347546 707162 348102 707718
rect 336986 698058 337542 698614
rect 336986 662058 337542 662614
rect 336986 626058 337542 626614
rect 336986 590058 337542 590614
rect 336986 554058 337542 554614
rect 336986 518058 337542 518614
rect 343826 705242 344382 705798
rect 343826 668898 344382 669454
rect 343826 632898 344382 633454
rect 343826 596898 344382 597454
rect 343826 560898 344382 561454
rect 343826 524898 344382 525454
rect 347546 672618 348102 673174
rect 347546 636618 348102 637174
rect 347546 600618 348102 601174
rect 347546 564618 348102 565174
rect 347546 528618 348102 529174
rect 347546 492618 348102 493174
rect 351266 676338 351822 676894
rect 351266 640338 351822 640894
rect 351266 604338 351822 604894
rect 351266 568338 351822 568894
rect 351266 532338 351822 532894
rect 351266 496338 351822 496894
rect 372986 710042 373542 710598
rect 369266 708122 369822 708678
rect 365546 706202 366102 706758
rect 354986 680058 355542 680614
rect 354986 644058 355542 644614
rect 354986 608058 355542 608614
rect 354986 572058 355542 572614
rect 354986 536058 355542 536614
rect 354986 500058 355542 500614
rect 361826 704282 362382 704838
rect 361826 686898 362382 687454
rect 361826 650898 362382 651454
rect 361826 614898 362382 615454
rect 361826 578898 362382 579454
rect 361826 542898 362382 543454
rect 361826 506898 362382 507454
rect 365546 690618 366102 691174
rect 365546 654618 366102 655174
rect 365546 618618 366102 619174
rect 365546 582618 366102 583174
rect 365546 546618 366102 547174
rect 365546 510618 366102 511174
rect 369266 694338 369822 694894
rect 369266 658338 369822 658894
rect 369266 622338 369822 622894
rect 369266 586338 369822 586894
rect 369266 550338 369822 550894
rect 369266 514338 369822 514894
rect 390986 711002 391542 711558
rect 387266 709082 387822 709638
rect 383546 707162 384102 707718
rect 372986 698058 373542 698614
rect 372986 662058 373542 662614
rect 372986 626058 373542 626614
rect 372986 590058 373542 590614
rect 372986 554058 373542 554614
rect 372986 518058 373542 518614
rect 379826 705242 380382 705798
rect 379826 668898 380382 669454
rect 379826 632898 380382 633454
rect 379826 596898 380382 597454
rect 379826 560898 380382 561454
rect 379826 524898 380382 525454
rect 383546 672618 384102 673174
rect 383546 636618 384102 637174
rect 383546 600618 384102 601174
rect 383546 564618 384102 565174
rect 383546 528618 384102 529174
rect 383546 492618 384102 493174
rect 387266 676338 387822 676894
rect 387266 640338 387822 640894
rect 387266 604338 387822 604894
rect 387266 568338 387822 568894
rect 387266 532338 387822 532894
rect 387266 496338 387822 496894
rect 228986 482058 229542 482614
rect 239250 471218 239486 471454
rect 239250 470898 239486 471134
rect 269970 471218 270206 471454
rect 269970 470898 270206 471134
rect 300690 471218 300926 471454
rect 300690 470898 300926 471134
rect 331410 471218 331646 471454
rect 331410 470898 331646 471134
rect 362130 471218 362366 471454
rect 362130 470898 362366 471134
rect 387266 460338 387822 460894
rect 254610 453218 254846 453454
rect 254610 452898 254846 453134
rect 285330 453218 285566 453454
rect 285330 452898 285566 453134
rect 316050 453218 316286 453454
rect 316050 452898 316286 453134
rect 346770 453218 347006 453454
rect 346770 452898 347006 453134
rect 377490 453218 377726 453454
rect 377490 452898 377726 453134
rect 228986 446058 229542 446614
rect 239250 435218 239486 435454
rect 239250 434898 239486 435134
rect 269970 435218 270206 435454
rect 269970 434898 270206 435134
rect 300690 435218 300926 435454
rect 300690 434898 300926 435134
rect 331410 435218 331646 435454
rect 331410 434898 331646 435134
rect 362130 435218 362366 435454
rect 362130 434898 362366 435134
rect 387266 424338 387822 424894
rect 254610 417218 254846 417454
rect 254610 416898 254846 417134
rect 285330 417218 285566 417454
rect 285330 416898 285566 417134
rect 316050 417218 316286 417454
rect 316050 416898 316286 417134
rect 346770 417218 347006 417454
rect 346770 416898 347006 417134
rect 377490 417218 377726 417454
rect 377490 416898 377726 417134
rect 228986 410058 229542 410614
rect 239250 399218 239486 399454
rect 239250 398898 239486 399134
rect 269970 399218 270206 399454
rect 269970 398898 270206 399134
rect 300690 399218 300926 399454
rect 300690 398898 300926 399134
rect 331410 399218 331646 399454
rect 331410 398898 331646 399134
rect 362130 399218 362366 399454
rect 362130 398898 362366 399134
rect 387266 388338 387822 388894
rect 254610 381218 254846 381454
rect 254610 380898 254846 381134
rect 285330 381218 285566 381454
rect 285330 380898 285566 381134
rect 316050 381218 316286 381454
rect 316050 380898 316286 381134
rect 346770 381218 347006 381454
rect 346770 380898 347006 381134
rect 377490 381218 377726 381454
rect 377490 380898 377726 381134
rect 228986 374058 229542 374614
rect 239250 363218 239486 363454
rect 239250 362898 239486 363134
rect 269970 363218 270206 363454
rect 269970 362898 270206 363134
rect 300690 363218 300926 363454
rect 300690 362898 300926 363134
rect 331410 363218 331646 363454
rect 331410 362898 331646 363134
rect 362130 363218 362366 363454
rect 362130 362898 362366 363134
rect 387266 352338 387822 352894
rect 254610 345218 254846 345454
rect 254610 344898 254846 345134
rect 285330 345218 285566 345454
rect 285330 344898 285566 345134
rect 316050 345218 316286 345454
rect 316050 344898 316286 345134
rect 346770 345218 347006 345454
rect 346770 344898 347006 345134
rect 377490 345218 377726 345454
rect 377490 344898 377726 345134
rect 228986 338058 229542 338614
rect 228986 302058 229542 302614
rect 228986 266058 229542 266614
rect 228986 230058 229542 230614
rect 228986 194058 229542 194614
rect 228986 158058 229542 158614
rect 228986 122058 229542 122614
rect 228986 86058 229542 86614
rect 228986 50058 229542 50614
rect 228986 14058 229542 14614
rect 210986 -7622 211542 -7066
rect 235826 308898 236382 309454
rect 235826 272898 236382 273454
rect 235826 236898 236382 237454
rect 235826 200898 236382 201454
rect 235826 164898 236382 165454
rect 235826 128898 236382 129454
rect 235826 92898 236382 93454
rect 235826 56898 236382 57454
rect 235826 20898 236382 21454
rect 235826 -1862 236382 -1306
rect 239546 312618 240102 313174
rect 239546 276618 240102 277174
rect 239546 240618 240102 241174
rect 239546 204618 240102 205174
rect 239546 168618 240102 169174
rect 239546 132618 240102 133174
rect 239546 96618 240102 97174
rect 239546 60618 240102 61174
rect 239546 24618 240102 25174
rect 239546 -3782 240102 -3226
rect 243266 316338 243822 316894
rect 243266 280338 243822 280894
rect 243266 244338 243822 244894
rect 243266 208338 243822 208894
rect 243266 172338 243822 172894
rect 243266 136338 243822 136894
rect 243266 100338 243822 100894
rect 243266 64338 243822 64894
rect 243266 28338 243822 28894
rect 243266 -5702 243822 -5146
rect 246986 320058 247542 320614
rect 246986 284058 247542 284614
rect 246986 248058 247542 248614
rect 246986 212058 247542 212614
rect 246986 176058 247542 176614
rect 246986 140058 247542 140614
rect 246986 104058 247542 104614
rect 246986 68058 247542 68614
rect 246986 32058 247542 32614
rect 228986 -6662 229542 -6106
rect 253826 326898 254382 327454
rect 253826 290898 254382 291454
rect 253826 254898 254382 255454
rect 253826 218898 254382 219454
rect 253826 182898 254382 183454
rect 253826 146898 254382 147454
rect 253826 110898 254382 111454
rect 253826 74898 254382 75454
rect 253826 38898 254382 39454
rect 253826 2898 254382 3454
rect 253826 -902 254382 -346
rect 257546 330618 258102 331174
rect 257546 294618 258102 295174
rect 257546 258618 258102 259174
rect 257546 222618 258102 223174
rect 257546 186618 258102 187174
rect 257546 150618 258102 151174
rect 257546 114618 258102 115174
rect 257546 78618 258102 79174
rect 257546 42618 258102 43174
rect 257546 6618 258102 7174
rect 257546 -2822 258102 -2266
rect 261266 334338 261822 334894
rect 261266 298338 261822 298894
rect 261266 262338 261822 262894
rect 261266 226338 261822 226894
rect 261266 190338 261822 190894
rect 261266 154338 261822 154894
rect 261266 118338 261822 118894
rect 261266 82338 261822 82894
rect 261266 46338 261822 46894
rect 261266 10338 261822 10894
rect 261266 -4742 261822 -4186
rect 264986 302058 265542 302614
rect 264986 266058 265542 266614
rect 264986 230058 265542 230614
rect 264986 194058 265542 194614
rect 264986 158058 265542 158614
rect 264986 122058 265542 122614
rect 264986 86058 265542 86614
rect 264986 50058 265542 50614
rect 264986 14058 265542 14614
rect 246986 -7622 247542 -7066
rect 271826 308898 272382 309454
rect 271826 272898 272382 273454
rect 271826 236898 272382 237454
rect 271826 200898 272382 201454
rect 271826 164898 272382 165454
rect 271826 128898 272382 129454
rect 271826 92898 272382 93454
rect 271826 56898 272382 57454
rect 271826 20898 272382 21454
rect 271826 -1862 272382 -1306
rect 275546 312618 276102 313174
rect 275546 276618 276102 277174
rect 275546 240618 276102 241174
rect 275546 204618 276102 205174
rect 275546 168618 276102 169174
rect 275546 132618 276102 133174
rect 275546 96618 276102 97174
rect 275546 60618 276102 61174
rect 275546 24618 276102 25174
rect 275546 -3782 276102 -3226
rect 279266 316338 279822 316894
rect 279266 280338 279822 280894
rect 279266 244338 279822 244894
rect 279266 208338 279822 208894
rect 279266 172338 279822 172894
rect 279266 136338 279822 136894
rect 279266 100338 279822 100894
rect 279266 64338 279822 64894
rect 279266 28338 279822 28894
rect 279266 -5702 279822 -5146
rect 282986 320058 283542 320614
rect 282986 284058 283542 284614
rect 282986 248058 283542 248614
rect 282986 212058 283542 212614
rect 282986 176058 283542 176614
rect 282986 140058 283542 140614
rect 282986 104058 283542 104614
rect 282986 68058 283542 68614
rect 282986 32058 283542 32614
rect 264986 -6662 265542 -6106
rect 289826 326898 290382 327454
rect 289826 290898 290382 291454
rect 289826 254898 290382 255454
rect 289826 218898 290382 219454
rect 289826 182898 290382 183454
rect 289826 146898 290382 147454
rect 289826 110898 290382 111454
rect 289826 74898 290382 75454
rect 289826 38898 290382 39454
rect 289826 2898 290382 3454
rect 289826 -902 290382 -346
rect 293546 330618 294102 331174
rect 293546 294618 294102 295174
rect 293546 258618 294102 259174
rect 293546 222618 294102 223174
rect 293546 186618 294102 187174
rect 293546 150618 294102 151174
rect 293546 114618 294102 115174
rect 293546 78618 294102 79174
rect 293546 42618 294102 43174
rect 293546 6618 294102 7174
rect 293546 -2822 294102 -2266
rect 297266 334338 297822 334894
rect 297266 298338 297822 298894
rect 297266 262338 297822 262894
rect 297266 226338 297822 226894
rect 297266 190338 297822 190894
rect 297266 154338 297822 154894
rect 297266 118338 297822 118894
rect 297266 82338 297822 82894
rect 297266 46338 297822 46894
rect 297266 10338 297822 10894
rect 297266 -4742 297822 -4186
rect 300986 302058 301542 302614
rect 300986 266058 301542 266614
rect 300986 230058 301542 230614
rect 300986 194058 301542 194614
rect 300986 158058 301542 158614
rect 300986 122058 301542 122614
rect 300986 86058 301542 86614
rect 300986 50058 301542 50614
rect 300986 14058 301542 14614
rect 282986 -7622 283542 -7066
rect 307826 308898 308382 309454
rect 307826 272898 308382 273454
rect 307826 236898 308382 237454
rect 307826 200898 308382 201454
rect 307826 164898 308382 165454
rect 307826 128898 308382 129454
rect 307826 92898 308382 93454
rect 307826 56898 308382 57454
rect 307826 20898 308382 21454
rect 307826 -1862 308382 -1306
rect 311546 312618 312102 313174
rect 311546 276618 312102 277174
rect 311546 240618 312102 241174
rect 311546 204618 312102 205174
rect 311546 168618 312102 169174
rect 311546 132618 312102 133174
rect 311546 96618 312102 97174
rect 311546 60618 312102 61174
rect 311546 24618 312102 25174
rect 311546 -3782 312102 -3226
rect 315266 316338 315822 316894
rect 315266 280338 315822 280894
rect 315266 244338 315822 244894
rect 315266 208338 315822 208894
rect 315266 172338 315822 172894
rect 315266 136338 315822 136894
rect 315266 100338 315822 100894
rect 315266 64338 315822 64894
rect 315266 28338 315822 28894
rect 315266 -5702 315822 -5146
rect 318986 320058 319542 320614
rect 318986 284058 319542 284614
rect 318986 248058 319542 248614
rect 318986 212058 319542 212614
rect 318986 176058 319542 176614
rect 318986 140058 319542 140614
rect 318986 104058 319542 104614
rect 318986 68058 319542 68614
rect 318986 32058 319542 32614
rect 300986 -6662 301542 -6106
rect 325826 326898 326382 327454
rect 325826 290898 326382 291454
rect 325826 254898 326382 255454
rect 325826 218898 326382 219454
rect 325826 182898 326382 183454
rect 325826 146898 326382 147454
rect 325826 110898 326382 111454
rect 325826 74898 326382 75454
rect 325826 38898 326382 39454
rect 325826 2898 326382 3454
rect 325826 -902 326382 -346
rect 329546 330618 330102 331174
rect 329546 294618 330102 295174
rect 329546 258618 330102 259174
rect 329546 222618 330102 223174
rect 329546 186618 330102 187174
rect 329546 150618 330102 151174
rect 329546 114618 330102 115174
rect 329546 78618 330102 79174
rect 329546 42618 330102 43174
rect 329546 6618 330102 7174
rect 329546 -2822 330102 -2266
rect 333266 334338 333822 334894
rect 333266 298338 333822 298894
rect 333266 262338 333822 262894
rect 333266 226338 333822 226894
rect 333266 190338 333822 190894
rect 333266 154338 333822 154894
rect 333266 118338 333822 118894
rect 333266 82338 333822 82894
rect 333266 46338 333822 46894
rect 333266 10338 333822 10894
rect 333266 -4742 333822 -4186
rect 336986 302058 337542 302614
rect 336986 266058 337542 266614
rect 336986 230058 337542 230614
rect 336986 194058 337542 194614
rect 336986 158058 337542 158614
rect 336986 122058 337542 122614
rect 336986 86058 337542 86614
rect 336986 50058 337542 50614
rect 336986 14058 337542 14614
rect 318986 -7622 319542 -7066
rect 343826 308898 344382 309454
rect 343826 272898 344382 273454
rect 343826 236898 344382 237454
rect 343826 200898 344382 201454
rect 343826 164898 344382 165454
rect 343826 128898 344382 129454
rect 343826 92898 344382 93454
rect 343826 56898 344382 57454
rect 343826 20898 344382 21454
rect 343826 -1862 344382 -1306
rect 347546 312618 348102 313174
rect 347546 276618 348102 277174
rect 347546 240618 348102 241174
rect 347546 204618 348102 205174
rect 347546 168618 348102 169174
rect 347546 132618 348102 133174
rect 347546 96618 348102 97174
rect 347546 60618 348102 61174
rect 347546 24618 348102 25174
rect 347546 -3782 348102 -3226
rect 351266 316338 351822 316894
rect 351266 280338 351822 280894
rect 351266 244338 351822 244894
rect 351266 208338 351822 208894
rect 351266 172338 351822 172894
rect 351266 136338 351822 136894
rect 351266 100338 351822 100894
rect 351266 64338 351822 64894
rect 351266 28338 351822 28894
rect 351266 -5702 351822 -5146
rect 354986 320058 355542 320614
rect 354986 284058 355542 284614
rect 354986 248058 355542 248614
rect 354986 212058 355542 212614
rect 354986 176058 355542 176614
rect 354986 140058 355542 140614
rect 354986 104058 355542 104614
rect 354986 68058 355542 68614
rect 354986 32058 355542 32614
rect 336986 -6662 337542 -6106
rect 361826 326898 362382 327454
rect 361826 290898 362382 291454
rect 361826 254898 362382 255454
rect 361826 218898 362382 219454
rect 361826 182898 362382 183454
rect 361826 146898 362382 147454
rect 361826 110898 362382 111454
rect 361826 74898 362382 75454
rect 361826 38898 362382 39454
rect 361826 2898 362382 3454
rect 361826 -902 362382 -346
rect 365546 330618 366102 331174
rect 365546 294618 366102 295174
rect 365546 258618 366102 259174
rect 365546 222618 366102 223174
rect 365546 186618 366102 187174
rect 365546 150618 366102 151174
rect 365546 114618 366102 115174
rect 365546 78618 366102 79174
rect 365546 42618 366102 43174
rect 365546 6618 366102 7174
rect 365546 -2822 366102 -2266
rect 369266 334338 369822 334894
rect 369266 298338 369822 298894
rect 369266 262338 369822 262894
rect 369266 226338 369822 226894
rect 369266 190338 369822 190894
rect 369266 154338 369822 154894
rect 369266 118338 369822 118894
rect 369266 82338 369822 82894
rect 369266 46338 369822 46894
rect 369266 10338 369822 10894
rect 369266 -4742 369822 -4186
rect 372986 302058 373542 302614
rect 372986 266058 373542 266614
rect 372986 230058 373542 230614
rect 372986 194058 373542 194614
rect 372986 158058 373542 158614
rect 372986 122058 373542 122614
rect 372986 86058 373542 86614
rect 372986 50058 373542 50614
rect 372986 14058 373542 14614
rect 354986 -7622 355542 -7066
rect 379826 308898 380382 309454
rect 379826 272898 380382 273454
rect 379826 236898 380382 237454
rect 379826 200898 380382 201454
rect 379826 164898 380382 165454
rect 379826 128898 380382 129454
rect 379826 92898 380382 93454
rect 379826 56898 380382 57454
rect 379826 20898 380382 21454
rect 379826 -1862 380382 -1306
rect 383546 312618 384102 313174
rect 383546 276618 384102 277174
rect 383546 240618 384102 241174
rect 383546 204618 384102 205174
rect 383546 168618 384102 169174
rect 383546 132618 384102 133174
rect 383546 96618 384102 97174
rect 383546 60618 384102 61174
rect 383546 24618 384102 25174
rect 383546 -3782 384102 -3226
rect 387266 316338 387822 316894
rect 387266 280338 387822 280894
rect 387266 244338 387822 244894
rect 387266 208338 387822 208894
rect 387266 172338 387822 172894
rect 387266 136338 387822 136894
rect 387266 100338 387822 100894
rect 387266 64338 387822 64894
rect 387266 28338 387822 28894
rect 387266 -5702 387822 -5146
rect 408986 710042 409542 710598
rect 405266 708122 405822 708678
rect 401546 706202 402102 706758
rect 390986 680058 391542 680614
rect 390986 644058 391542 644614
rect 390986 608058 391542 608614
rect 390986 572058 391542 572614
rect 390986 536058 391542 536614
rect 390986 500058 391542 500614
rect 390986 464058 391542 464614
rect 390986 428058 391542 428614
rect 390986 392058 391542 392614
rect 390986 356058 391542 356614
rect 390986 320058 391542 320614
rect 390986 284058 391542 284614
rect 390986 248058 391542 248614
rect 390986 212058 391542 212614
rect 390986 176058 391542 176614
rect 390986 140058 391542 140614
rect 390986 104058 391542 104614
rect 390986 68058 391542 68614
rect 390986 32058 391542 32614
rect 372986 -6662 373542 -6106
rect 397826 704282 398382 704838
rect 397826 686898 398382 687454
rect 397826 650898 398382 651454
rect 397826 614898 398382 615454
rect 397826 578898 398382 579454
rect 397826 542898 398382 543454
rect 397826 506898 398382 507454
rect 397826 470898 398382 471454
rect 397826 434898 398382 435454
rect 397826 398898 398382 399454
rect 397826 362898 398382 363454
rect 397826 326898 398382 327454
rect 397826 290898 398382 291454
rect 397826 254898 398382 255454
rect 397826 218898 398382 219454
rect 397826 182898 398382 183454
rect 397826 146898 398382 147454
rect 397826 110898 398382 111454
rect 397826 74898 398382 75454
rect 397826 38898 398382 39454
rect 397826 2898 398382 3454
rect 397826 -902 398382 -346
rect 401546 690618 402102 691174
rect 401546 654618 402102 655174
rect 401546 618618 402102 619174
rect 401546 582618 402102 583174
rect 401546 546618 402102 547174
rect 401546 510618 402102 511174
rect 401546 474618 402102 475174
rect 401546 438618 402102 439174
rect 401546 402618 402102 403174
rect 401546 366618 402102 367174
rect 401546 330618 402102 331174
rect 401546 294618 402102 295174
rect 401546 258618 402102 259174
rect 401546 222618 402102 223174
rect 401546 186618 402102 187174
rect 401546 150618 402102 151174
rect 401546 114618 402102 115174
rect 401546 78618 402102 79174
rect 401546 42618 402102 43174
rect 401546 6618 402102 7174
rect 401546 -2822 402102 -2266
rect 405266 694338 405822 694894
rect 405266 658338 405822 658894
rect 405266 622338 405822 622894
rect 405266 586338 405822 586894
rect 405266 550338 405822 550894
rect 405266 514338 405822 514894
rect 405266 478338 405822 478894
rect 405266 442338 405822 442894
rect 405266 406338 405822 406894
rect 405266 370338 405822 370894
rect 405266 334338 405822 334894
rect 405266 298338 405822 298894
rect 405266 262338 405822 262894
rect 405266 226338 405822 226894
rect 405266 190338 405822 190894
rect 405266 154338 405822 154894
rect 405266 118338 405822 118894
rect 405266 82338 405822 82894
rect 405266 46338 405822 46894
rect 405266 10338 405822 10894
rect 405266 -4742 405822 -4186
rect 426986 711002 427542 711558
rect 423266 709082 423822 709638
rect 419546 707162 420102 707718
rect 408986 698058 409542 698614
rect 408986 662058 409542 662614
rect 408986 626058 409542 626614
rect 408986 590058 409542 590614
rect 408986 554058 409542 554614
rect 408986 518058 409542 518614
rect 408986 482058 409542 482614
rect 408986 446058 409542 446614
rect 408986 410058 409542 410614
rect 408986 374058 409542 374614
rect 408986 338058 409542 338614
rect 408986 302058 409542 302614
rect 408986 266058 409542 266614
rect 408986 230058 409542 230614
rect 408986 194058 409542 194614
rect 408986 158058 409542 158614
rect 408986 122058 409542 122614
rect 408986 86058 409542 86614
rect 408986 50058 409542 50614
rect 408986 14058 409542 14614
rect 390986 -7622 391542 -7066
rect 415826 705242 416382 705798
rect 415826 668898 416382 669454
rect 415826 632898 416382 633454
rect 415826 596898 416382 597454
rect 415826 560898 416382 561454
rect 415826 524898 416382 525454
rect 415826 488898 416382 489454
rect 415826 452898 416382 453454
rect 415826 416898 416382 417454
rect 415826 380898 416382 381454
rect 415826 344898 416382 345454
rect 415826 308898 416382 309454
rect 415826 272898 416382 273454
rect 415826 236898 416382 237454
rect 415826 200898 416382 201454
rect 415826 164898 416382 165454
rect 415826 128898 416382 129454
rect 415826 92898 416382 93454
rect 415826 56898 416382 57454
rect 415826 20898 416382 21454
rect 415826 -1862 416382 -1306
rect 419546 672618 420102 673174
rect 419546 636618 420102 637174
rect 419546 600618 420102 601174
rect 419546 564618 420102 565174
rect 419546 528618 420102 529174
rect 419546 492618 420102 493174
rect 419546 456618 420102 457174
rect 419546 420618 420102 421174
rect 419546 384618 420102 385174
rect 419546 348618 420102 349174
rect 419546 312618 420102 313174
rect 419546 276618 420102 277174
rect 419546 240618 420102 241174
rect 419546 204618 420102 205174
rect 419546 168618 420102 169174
rect 419546 132618 420102 133174
rect 419546 96618 420102 97174
rect 419546 60618 420102 61174
rect 419546 24618 420102 25174
rect 419546 -3782 420102 -3226
rect 423266 676338 423822 676894
rect 423266 640338 423822 640894
rect 423266 604338 423822 604894
rect 423266 568338 423822 568894
rect 423266 532338 423822 532894
rect 423266 496338 423822 496894
rect 423266 460338 423822 460894
rect 423266 424338 423822 424894
rect 423266 388338 423822 388894
rect 423266 352338 423822 352894
rect 423266 316338 423822 316894
rect 423266 280338 423822 280894
rect 423266 244338 423822 244894
rect 423266 208338 423822 208894
rect 423266 172338 423822 172894
rect 423266 136338 423822 136894
rect 423266 100338 423822 100894
rect 423266 64338 423822 64894
rect 423266 28338 423822 28894
rect 423266 -5702 423822 -5146
rect 444986 710042 445542 710598
rect 441266 708122 441822 708678
rect 437546 706202 438102 706758
rect 426986 680058 427542 680614
rect 426986 644058 427542 644614
rect 426986 608058 427542 608614
rect 426986 572058 427542 572614
rect 426986 536058 427542 536614
rect 426986 500058 427542 500614
rect 426986 464058 427542 464614
rect 426986 428058 427542 428614
rect 426986 392058 427542 392614
rect 426986 356058 427542 356614
rect 426986 320058 427542 320614
rect 426986 284058 427542 284614
rect 426986 248058 427542 248614
rect 426986 212058 427542 212614
rect 426986 176058 427542 176614
rect 426986 140058 427542 140614
rect 426986 104058 427542 104614
rect 426986 68058 427542 68614
rect 426986 32058 427542 32614
rect 408986 -6662 409542 -6106
rect 433826 704282 434382 704838
rect 433826 686898 434382 687454
rect 433826 650898 434382 651454
rect 433826 614898 434382 615454
rect 433826 578898 434382 579454
rect 433826 542898 434382 543454
rect 433826 506898 434382 507454
rect 433826 470898 434382 471454
rect 433826 434898 434382 435454
rect 433826 398898 434382 399454
rect 433826 362898 434382 363454
rect 433826 326898 434382 327454
rect 433826 290898 434382 291454
rect 433826 254898 434382 255454
rect 433826 218898 434382 219454
rect 433826 182898 434382 183454
rect 433826 146898 434382 147454
rect 433826 110898 434382 111454
rect 433826 74898 434382 75454
rect 433826 38898 434382 39454
rect 433826 2898 434382 3454
rect 433826 -902 434382 -346
rect 437546 690618 438102 691174
rect 437546 654618 438102 655174
rect 437546 618618 438102 619174
rect 437546 582618 438102 583174
rect 437546 546618 438102 547174
rect 437546 510618 438102 511174
rect 437546 474618 438102 475174
rect 437546 438618 438102 439174
rect 437546 402618 438102 403174
rect 437546 366618 438102 367174
rect 437546 330618 438102 331174
rect 437546 294618 438102 295174
rect 437546 258618 438102 259174
rect 437546 222618 438102 223174
rect 437546 186618 438102 187174
rect 437546 150618 438102 151174
rect 437546 114618 438102 115174
rect 437546 78618 438102 79174
rect 437546 42618 438102 43174
rect 437546 6618 438102 7174
rect 437546 -2822 438102 -2266
rect 441266 694338 441822 694894
rect 441266 658338 441822 658894
rect 441266 622338 441822 622894
rect 441266 586338 441822 586894
rect 441266 550338 441822 550894
rect 441266 514338 441822 514894
rect 441266 478338 441822 478894
rect 441266 442338 441822 442894
rect 441266 406338 441822 406894
rect 441266 370338 441822 370894
rect 441266 334338 441822 334894
rect 441266 298338 441822 298894
rect 441266 262338 441822 262894
rect 441266 226338 441822 226894
rect 441266 190338 441822 190894
rect 441266 154338 441822 154894
rect 441266 118338 441822 118894
rect 441266 82338 441822 82894
rect 441266 46338 441822 46894
rect 441266 10338 441822 10894
rect 441266 -4742 441822 -4186
rect 462986 711002 463542 711558
rect 459266 709082 459822 709638
rect 455546 707162 456102 707718
rect 444986 698058 445542 698614
rect 444986 662058 445542 662614
rect 444986 626058 445542 626614
rect 444986 590058 445542 590614
rect 444986 554058 445542 554614
rect 444986 518058 445542 518614
rect 444986 482058 445542 482614
rect 444986 446058 445542 446614
rect 444986 410058 445542 410614
rect 444986 374058 445542 374614
rect 444986 338058 445542 338614
rect 444986 302058 445542 302614
rect 444986 266058 445542 266614
rect 444986 230058 445542 230614
rect 444986 194058 445542 194614
rect 444986 158058 445542 158614
rect 444986 122058 445542 122614
rect 444986 86058 445542 86614
rect 444986 50058 445542 50614
rect 444986 14058 445542 14614
rect 426986 -7622 427542 -7066
rect 451826 705242 452382 705798
rect 451826 668898 452382 669454
rect 451826 632898 452382 633454
rect 451826 596898 452382 597454
rect 451826 560898 452382 561454
rect 451826 524898 452382 525454
rect 451826 488898 452382 489454
rect 451826 452898 452382 453454
rect 451826 416898 452382 417454
rect 451826 380898 452382 381454
rect 451826 344898 452382 345454
rect 451826 308898 452382 309454
rect 451826 272898 452382 273454
rect 451826 236898 452382 237454
rect 451826 200898 452382 201454
rect 451826 164898 452382 165454
rect 451826 128898 452382 129454
rect 451826 92898 452382 93454
rect 451826 56898 452382 57454
rect 451826 20898 452382 21454
rect 451826 -1862 452382 -1306
rect 455546 672618 456102 673174
rect 455546 636618 456102 637174
rect 455546 600618 456102 601174
rect 455546 564618 456102 565174
rect 455546 528618 456102 529174
rect 455546 492618 456102 493174
rect 455546 456618 456102 457174
rect 455546 420618 456102 421174
rect 455546 384618 456102 385174
rect 455546 348618 456102 349174
rect 455546 312618 456102 313174
rect 455546 276618 456102 277174
rect 455546 240618 456102 241174
rect 455546 204618 456102 205174
rect 455546 168618 456102 169174
rect 455546 132618 456102 133174
rect 455546 96618 456102 97174
rect 455546 60618 456102 61174
rect 455546 24618 456102 25174
rect 455546 -3782 456102 -3226
rect 459266 676338 459822 676894
rect 459266 640338 459822 640894
rect 459266 604338 459822 604894
rect 459266 568338 459822 568894
rect 459266 532338 459822 532894
rect 459266 496338 459822 496894
rect 459266 460338 459822 460894
rect 459266 424338 459822 424894
rect 459266 388338 459822 388894
rect 459266 352338 459822 352894
rect 459266 316338 459822 316894
rect 459266 280338 459822 280894
rect 459266 244338 459822 244894
rect 459266 208338 459822 208894
rect 459266 172338 459822 172894
rect 459266 136338 459822 136894
rect 459266 100338 459822 100894
rect 459266 64338 459822 64894
rect 459266 28338 459822 28894
rect 459266 -5702 459822 -5146
rect 480986 710042 481542 710598
rect 477266 708122 477822 708678
rect 473546 706202 474102 706758
rect 462986 680058 463542 680614
rect 462986 644058 463542 644614
rect 462986 608058 463542 608614
rect 462986 572058 463542 572614
rect 462986 536058 463542 536614
rect 462986 500058 463542 500614
rect 462986 464058 463542 464614
rect 462986 428058 463542 428614
rect 462986 392058 463542 392614
rect 462986 356058 463542 356614
rect 462986 320058 463542 320614
rect 462986 284058 463542 284614
rect 462986 248058 463542 248614
rect 462986 212058 463542 212614
rect 462986 176058 463542 176614
rect 462986 140058 463542 140614
rect 462986 104058 463542 104614
rect 462986 68058 463542 68614
rect 462986 32058 463542 32614
rect 444986 -6662 445542 -6106
rect 469826 704282 470382 704838
rect 469826 686898 470382 687454
rect 469826 650898 470382 651454
rect 469826 614898 470382 615454
rect 469826 578898 470382 579454
rect 469826 542898 470382 543454
rect 469826 506898 470382 507454
rect 469826 470898 470382 471454
rect 469826 434898 470382 435454
rect 469826 398898 470382 399454
rect 469826 362898 470382 363454
rect 469826 326898 470382 327454
rect 469826 290898 470382 291454
rect 469826 254898 470382 255454
rect 469826 218898 470382 219454
rect 469826 182898 470382 183454
rect 469826 146898 470382 147454
rect 469826 110898 470382 111454
rect 469826 74898 470382 75454
rect 469826 38898 470382 39454
rect 469826 2898 470382 3454
rect 469826 -902 470382 -346
rect 473546 690618 474102 691174
rect 473546 654618 474102 655174
rect 473546 618618 474102 619174
rect 473546 582618 474102 583174
rect 473546 546618 474102 547174
rect 473546 510618 474102 511174
rect 473546 474618 474102 475174
rect 473546 438618 474102 439174
rect 473546 402618 474102 403174
rect 473546 366618 474102 367174
rect 473546 330618 474102 331174
rect 473546 294618 474102 295174
rect 473546 258618 474102 259174
rect 473546 222618 474102 223174
rect 473546 186618 474102 187174
rect 473546 150618 474102 151174
rect 473546 114618 474102 115174
rect 473546 78618 474102 79174
rect 473546 42618 474102 43174
rect 473546 6618 474102 7174
rect 473546 -2822 474102 -2266
rect 477266 694338 477822 694894
rect 477266 658338 477822 658894
rect 477266 622338 477822 622894
rect 477266 586338 477822 586894
rect 477266 550338 477822 550894
rect 477266 514338 477822 514894
rect 477266 478338 477822 478894
rect 477266 442338 477822 442894
rect 477266 406338 477822 406894
rect 477266 370338 477822 370894
rect 477266 334338 477822 334894
rect 477266 298338 477822 298894
rect 477266 262338 477822 262894
rect 477266 226338 477822 226894
rect 477266 190338 477822 190894
rect 477266 154338 477822 154894
rect 477266 118338 477822 118894
rect 477266 82338 477822 82894
rect 477266 46338 477822 46894
rect 477266 10338 477822 10894
rect 477266 -4742 477822 -4186
rect 498986 711002 499542 711558
rect 495266 709082 495822 709638
rect 491546 707162 492102 707718
rect 480986 698058 481542 698614
rect 480986 662058 481542 662614
rect 480986 626058 481542 626614
rect 480986 590058 481542 590614
rect 480986 554058 481542 554614
rect 480986 518058 481542 518614
rect 480986 482058 481542 482614
rect 480986 446058 481542 446614
rect 480986 410058 481542 410614
rect 480986 374058 481542 374614
rect 480986 338058 481542 338614
rect 480986 302058 481542 302614
rect 480986 266058 481542 266614
rect 480986 230058 481542 230614
rect 480986 194058 481542 194614
rect 480986 158058 481542 158614
rect 480986 122058 481542 122614
rect 480986 86058 481542 86614
rect 480986 50058 481542 50614
rect 480986 14058 481542 14614
rect 462986 -7622 463542 -7066
rect 487826 705242 488382 705798
rect 487826 668898 488382 669454
rect 487826 632898 488382 633454
rect 487826 596898 488382 597454
rect 487826 560898 488382 561454
rect 487826 524898 488382 525454
rect 487826 488898 488382 489454
rect 487826 452898 488382 453454
rect 487826 416898 488382 417454
rect 487826 380898 488382 381454
rect 487826 344898 488382 345454
rect 487826 308898 488382 309454
rect 487826 272898 488382 273454
rect 487826 236898 488382 237454
rect 487826 200898 488382 201454
rect 487826 164898 488382 165454
rect 487826 128898 488382 129454
rect 487826 92898 488382 93454
rect 487826 56898 488382 57454
rect 487826 20898 488382 21454
rect 487826 -1862 488382 -1306
rect 491546 672618 492102 673174
rect 491546 636618 492102 637174
rect 491546 600618 492102 601174
rect 491546 564618 492102 565174
rect 491546 528618 492102 529174
rect 491546 492618 492102 493174
rect 491546 456618 492102 457174
rect 491546 420618 492102 421174
rect 491546 384618 492102 385174
rect 491546 348618 492102 349174
rect 491546 312618 492102 313174
rect 491546 276618 492102 277174
rect 491546 240618 492102 241174
rect 491546 204618 492102 205174
rect 491546 168618 492102 169174
rect 491546 132618 492102 133174
rect 491546 96618 492102 97174
rect 491546 60618 492102 61174
rect 491546 24618 492102 25174
rect 491546 -3782 492102 -3226
rect 495266 676338 495822 676894
rect 495266 640338 495822 640894
rect 495266 604338 495822 604894
rect 495266 568338 495822 568894
rect 495266 532338 495822 532894
rect 495266 496338 495822 496894
rect 495266 460338 495822 460894
rect 495266 424338 495822 424894
rect 495266 388338 495822 388894
rect 495266 352338 495822 352894
rect 495266 316338 495822 316894
rect 495266 280338 495822 280894
rect 495266 244338 495822 244894
rect 495266 208338 495822 208894
rect 495266 172338 495822 172894
rect 495266 136338 495822 136894
rect 495266 100338 495822 100894
rect 495266 64338 495822 64894
rect 495266 28338 495822 28894
rect 495266 -5702 495822 -5146
rect 516986 710042 517542 710598
rect 513266 708122 513822 708678
rect 509546 706202 510102 706758
rect 498986 680058 499542 680614
rect 498986 644058 499542 644614
rect 498986 608058 499542 608614
rect 498986 572058 499542 572614
rect 498986 536058 499542 536614
rect 498986 500058 499542 500614
rect 498986 464058 499542 464614
rect 498986 428058 499542 428614
rect 498986 392058 499542 392614
rect 498986 356058 499542 356614
rect 498986 320058 499542 320614
rect 498986 284058 499542 284614
rect 498986 248058 499542 248614
rect 498986 212058 499542 212614
rect 498986 176058 499542 176614
rect 498986 140058 499542 140614
rect 498986 104058 499542 104614
rect 498986 68058 499542 68614
rect 498986 32058 499542 32614
rect 480986 -6662 481542 -6106
rect 505826 704282 506382 704838
rect 505826 686898 506382 687454
rect 505826 650898 506382 651454
rect 505826 614898 506382 615454
rect 505826 578898 506382 579454
rect 505826 542898 506382 543454
rect 505826 506898 506382 507454
rect 505826 470898 506382 471454
rect 505826 434898 506382 435454
rect 505826 398898 506382 399454
rect 505826 362898 506382 363454
rect 505826 326898 506382 327454
rect 505826 290898 506382 291454
rect 505826 254898 506382 255454
rect 505826 218898 506382 219454
rect 505826 182898 506382 183454
rect 505826 146898 506382 147454
rect 505826 110898 506382 111454
rect 505826 74898 506382 75454
rect 505826 38898 506382 39454
rect 505826 2898 506382 3454
rect 505826 -902 506382 -346
rect 509546 690618 510102 691174
rect 509546 654618 510102 655174
rect 509546 618618 510102 619174
rect 509546 582618 510102 583174
rect 509546 546618 510102 547174
rect 509546 510618 510102 511174
rect 509546 474618 510102 475174
rect 509546 438618 510102 439174
rect 509546 402618 510102 403174
rect 509546 366618 510102 367174
rect 509546 330618 510102 331174
rect 509546 294618 510102 295174
rect 509546 258618 510102 259174
rect 509546 222618 510102 223174
rect 509546 186618 510102 187174
rect 509546 150618 510102 151174
rect 509546 114618 510102 115174
rect 509546 78618 510102 79174
rect 509546 42618 510102 43174
rect 509546 6618 510102 7174
rect 509546 -2822 510102 -2266
rect 513266 694338 513822 694894
rect 513266 658338 513822 658894
rect 513266 622338 513822 622894
rect 513266 586338 513822 586894
rect 513266 550338 513822 550894
rect 513266 514338 513822 514894
rect 513266 478338 513822 478894
rect 513266 442338 513822 442894
rect 513266 406338 513822 406894
rect 513266 370338 513822 370894
rect 513266 334338 513822 334894
rect 513266 298338 513822 298894
rect 513266 262338 513822 262894
rect 513266 226338 513822 226894
rect 513266 190338 513822 190894
rect 513266 154338 513822 154894
rect 513266 118338 513822 118894
rect 513266 82338 513822 82894
rect 513266 46338 513822 46894
rect 513266 10338 513822 10894
rect 513266 -4742 513822 -4186
rect 534986 711002 535542 711558
rect 531266 709082 531822 709638
rect 527546 707162 528102 707718
rect 516986 698058 517542 698614
rect 516986 662058 517542 662614
rect 516986 626058 517542 626614
rect 516986 590058 517542 590614
rect 516986 554058 517542 554614
rect 516986 518058 517542 518614
rect 516986 482058 517542 482614
rect 516986 446058 517542 446614
rect 516986 410058 517542 410614
rect 516986 374058 517542 374614
rect 516986 338058 517542 338614
rect 516986 302058 517542 302614
rect 516986 266058 517542 266614
rect 516986 230058 517542 230614
rect 516986 194058 517542 194614
rect 516986 158058 517542 158614
rect 516986 122058 517542 122614
rect 516986 86058 517542 86614
rect 516986 50058 517542 50614
rect 516986 14058 517542 14614
rect 498986 -7622 499542 -7066
rect 523826 705242 524382 705798
rect 523826 668898 524382 669454
rect 523826 632898 524382 633454
rect 523826 596898 524382 597454
rect 523826 560898 524382 561454
rect 523826 524898 524382 525454
rect 523826 488898 524382 489454
rect 523826 452898 524382 453454
rect 523826 416898 524382 417454
rect 523826 380898 524382 381454
rect 523826 344898 524382 345454
rect 523826 308898 524382 309454
rect 523826 272898 524382 273454
rect 523826 236898 524382 237454
rect 523826 200898 524382 201454
rect 523826 164898 524382 165454
rect 523826 128898 524382 129454
rect 523826 92898 524382 93454
rect 523826 56898 524382 57454
rect 523826 20898 524382 21454
rect 523826 -1862 524382 -1306
rect 527546 672618 528102 673174
rect 527546 636618 528102 637174
rect 527546 600618 528102 601174
rect 527546 564618 528102 565174
rect 527546 528618 528102 529174
rect 527546 492618 528102 493174
rect 527546 456618 528102 457174
rect 527546 420618 528102 421174
rect 527546 384618 528102 385174
rect 527546 348618 528102 349174
rect 527546 312618 528102 313174
rect 527546 276618 528102 277174
rect 527546 240618 528102 241174
rect 527546 204618 528102 205174
rect 527546 168618 528102 169174
rect 527546 132618 528102 133174
rect 527546 96618 528102 97174
rect 527546 60618 528102 61174
rect 527546 24618 528102 25174
rect 527546 -3782 528102 -3226
rect 531266 676338 531822 676894
rect 531266 640338 531822 640894
rect 531266 604338 531822 604894
rect 531266 568338 531822 568894
rect 531266 532338 531822 532894
rect 531266 496338 531822 496894
rect 531266 460338 531822 460894
rect 531266 424338 531822 424894
rect 531266 388338 531822 388894
rect 531266 352338 531822 352894
rect 531266 316338 531822 316894
rect 531266 280338 531822 280894
rect 531266 244338 531822 244894
rect 531266 208338 531822 208894
rect 531266 172338 531822 172894
rect 531266 136338 531822 136894
rect 531266 100338 531822 100894
rect 531266 64338 531822 64894
rect 531266 28338 531822 28894
rect 531266 -5702 531822 -5146
rect 552986 710042 553542 710598
rect 549266 708122 549822 708678
rect 545546 706202 546102 706758
rect 534986 680058 535542 680614
rect 534986 644058 535542 644614
rect 534986 608058 535542 608614
rect 534986 572058 535542 572614
rect 534986 536058 535542 536614
rect 534986 500058 535542 500614
rect 534986 464058 535542 464614
rect 534986 428058 535542 428614
rect 534986 392058 535542 392614
rect 534986 356058 535542 356614
rect 534986 320058 535542 320614
rect 534986 284058 535542 284614
rect 534986 248058 535542 248614
rect 534986 212058 535542 212614
rect 534986 176058 535542 176614
rect 534986 140058 535542 140614
rect 534986 104058 535542 104614
rect 534986 68058 535542 68614
rect 534986 32058 535542 32614
rect 516986 -6662 517542 -6106
rect 541826 704282 542382 704838
rect 541826 686898 542382 687454
rect 541826 650898 542382 651454
rect 541826 614898 542382 615454
rect 541826 578898 542382 579454
rect 541826 542898 542382 543454
rect 541826 506898 542382 507454
rect 541826 470898 542382 471454
rect 541826 434898 542382 435454
rect 541826 398898 542382 399454
rect 541826 362898 542382 363454
rect 541826 326898 542382 327454
rect 541826 290898 542382 291454
rect 541826 254898 542382 255454
rect 541826 218898 542382 219454
rect 541826 182898 542382 183454
rect 541826 146898 542382 147454
rect 541826 110898 542382 111454
rect 541826 74898 542382 75454
rect 541826 38898 542382 39454
rect 541826 2898 542382 3454
rect 541826 -902 542382 -346
rect 545546 690618 546102 691174
rect 545546 654618 546102 655174
rect 545546 618618 546102 619174
rect 545546 582618 546102 583174
rect 545546 546618 546102 547174
rect 545546 510618 546102 511174
rect 545546 474618 546102 475174
rect 545546 438618 546102 439174
rect 545546 402618 546102 403174
rect 545546 366618 546102 367174
rect 545546 330618 546102 331174
rect 545546 294618 546102 295174
rect 545546 258618 546102 259174
rect 545546 222618 546102 223174
rect 545546 186618 546102 187174
rect 545546 150618 546102 151174
rect 545546 114618 546102 115174
rect 545546 78618 546102 79174
rect 545546 42618 546102 43174
rect 545546 6618 546102 7174
rect 545546 -2822 546102 -2266
rect 549266 694338 549822 694894
rect 549266 658338 549822 658894
rect 549266 622338 549822 622894
rect 549266 586338 549822 586894
rect 549266 550338 549822 550894
rect 549266 514338 549822 514894
rect 549266 478338 549822 478894
rect 549266 442338 549822 442894
rect 549266 406338 549822 406894
rect 549266 370338 549822 370894
rect 549266 334338 549822 334894
rect 549266 298338 549822 298894
rect 549266 262338 549822 262894
rect 549266 226338 549822 226894
rect 549266 190338 549822 190894
rect 549266 154338 549822 154894
rect 549266 118338 549822 118894
rect 549266 82338 549822 82894
rect 549266 46338 549822 46894
rect 549266 10338 549822 10894
rect 549266 -4742 549822 -4186
rect 570986 711002 571542 711558
rect 567266 709082 567822 709638
rect 563546 707162 564102 707718
rect 552986 698058 553542 698614
rect 552986 662058 553542 662614
rect 552986 626058 553542 626614
rect 552986 590058 553542 590614
rect 552986 554058 553542 554614
rect 552986 518058 553542 518614
rect 552986 482058 553542 482614
rect 552986 446058 553542 446614
rect 552986 410058 553542 410614
rect 552986 374058 553542 374614
rect 552986 338058 553542 338614
rect 552986 302058 553542 302614
rect 552986 266058 553542 266614
rect 552986 230058 553542 230614
rect 552986 194058 553542 194614
rect 552986 158058 553542 158614
rect 552986 122058 553542 122614
rect 552986 86058 553542 86614
rect 552986 50058 553542 50614
rect 552986 14058 553542 14614
rect 534986 -7622 535542 -7066
rect 559826 705242 560382 705798
rect 559826 668898 560382 669454
rect 559826 632898 560382 633454
rect 559826 596898 560382 597454
rect 559826 560898 560382 561454
rect 559826 524898 560382 525454
rect 559826 488898 560382 489454
rect 559826 452898 560382 453454
rect 559826 416898 560382 417454
rect 559826 380898 560382 381454
rect 559826 344898 560382 345454
rect 559826 308898 560382 309454
rect 559826 272898 560382 273454
rect 559826 236898 560382 237454
rect 559826 200898 560382 201454
rect 559826 164898 560382 165454
rect 559826 128898 560382 129454
rect 559826 92898 560382 93454
rect 559826 56898 560382 57454
rect 559826 20898 560382 21454
rect 559826 -1862 560382 -1306
rect 563546 672618 564102 673174
rect 563546 636618 564102 637174
rect 563546 600618 564102 601174
rect 563546 564618 564102 565174
rect 563546 528618 564102 529174
rect 563546 492618 564102 493174
rect 563546 456618 564102 457174
rect 563546 420618 564102 421174
rect 563546 384618 564102 385174
rect 563546 348618 564102 349174
rect 563546 312618 564102 313174
rect 563546 276618 564102 277174
rect 563546 240618 564102 241174
rect 563546 204618 564102 205174
rect 563546 168618 564102 169174
rect 563546 132618 564102 133174
rect 563546 96618 564102 97174
rect 563546 60618 564102 61174
rect 563546 24618 564102 25174
rect 563546 -3782 564102 -3226
rect 567266 676338 567822 676894
rect 567266 640338 567822 640894
rect 567266 604338 567822 604894
rect 567266 568338 567822 568894
rect 567266 532338 567822 532894
rect 567266 496338 567822 496894
rect 567266 460338 567822 460894
rect 567266 424338 567822 424894
rect 567266 388338 567822 388894
rect 567266 352338 567822 352894
rect 567266 316338 567822 316894
rect 567266 280338 567822 280894
rect 567266 244338 567822 244894
rect 567266 208338 567822 208894
rect 567266 172338 567822 172894
rect 567266 136338 567822 136894
rect 567266 100338 567822 100894
rect 567266 64338 567822 64894
rect 567266 28338 567822 28894
rect 567266 -5702 567822 -5146
rect 592062 711002 592618 711558
rect 591102 710042 591658 710598
rect 590142 709082 590698 709638
rect 589182 708122 589738 708678
rect 588222 707162 588778 707718
rect 581546 706202 582102 706758
rect 570986 680058 571542 680614
rect 570986 644058 571542 644614
rect 570986 608058 571542 608614
rect 570986 572058 571542 572614
rect 570986 536058 571542 536614
rect 570986 500058 571542 500614
rect 570986 464058 571542 464614
rect 570986 428058 571542 428614
rect 570986 392058 571542 392614
rect 570986 356058 571542 356614
rect 570986 320058 571542 320614
rect 570986 284058 571542 284614
rect 570986 248058 571542 248614
rect 570986 212058 571542 212614
rect 570986 176058 571542 176614
rect 570986 140058 571542 140614
rect 570986 104058 571542 104614
rect 570986 68058 571542 68614
rect 570986 32058 571542 32614
rect 552986 -6662 553542 -6106
rect 577826 704282 578382 704838
rect 577826 686898 578382 687454
rect 577826 650898 578382 651454
rect 577826 614898 578382 615454
rect 577826 578898 578382 579454
rect 577826 542898 578382 543454
rect 577826 506898 578382 507454
rect 577826 470898 578382 471454
rect 577826 434898 578382 435454
rect 577826 398898 578382 399454
rect 577826 362898 578382 363454
rect 577826 326898 578382 327454
rect 577826 290898 578382 291454
rect 577826 254898 578382 255454
rect 577826 218898 578382 219454
rect 577826 182898 578382 183454
rect 577826 146898 578382 147454
rect 577826 110898 578382 111454
rect 577826 74898 578382 75454
rect 577826 38898 578382 39454
rect 577826 2898 578382 3454
rect 577826 -902 578382 -346
rect 587262 706202 587818 706758
rect 586302 705242 586858 705798
rect 581546 690618 582102 691174
rect 581546 654618 582102 655174
rect 581546 618618 582102 619174
rect 581546 582618 582102 583174
rect 581546 546618 582102 547174
rect 581546 510618 582102 511174
rect 581546 474618 582102 475174
rect 581546 438618 582102 439174
rect 581546 402618 582102 403174
rect 581546 366618 582102 367174
rect 581546 330618 582102 331174
rect 581546 294618 582102 295174
rect 581546 258618 582102 259174
rect 581546 222618 582102 223174
rect 581546 186618 582102 187174
rect 581546 150618 582102 151174
rect 581546 114618 582102 115174
rect 581546 78618 582102 79174
rect 581546 42618 582102 43174
rect 581546 6618 582102 7174
rect 585342 704282 585898 704838
rect 585342 686898 585898 687454
rect 585342 650898 585898 651454
rect 585342 614898 585898 615454
rect 585342 578898 585898 579454
rect 585342 542898 585898 543454
rect 585342 506898 585898 507454
rect 585342 470898 585898 471454
rect 585342 434898 585898 435454
rect 585342 398898 585898 399454
rect 585342 362898 585898 363454
rect 585342 326898 585898 327454
rect 585342 290898 585898 291454
rect 585342 254898 585898 255454
rect 585342 218898 585898 219454
rect 585342 182898 585898 183454
rect 585342 146898 585898 147454
rect 585342 110898 585898 111454
rect 585342 74898 585898 75454
rect 585342 38898 585898 39454
rect 585342 2898 585898 3454
rect 585342 -902 585898 -346
rect 586302 668898 586858 669454
rect 586302 632898 586858 633454
rect 586302 596898 586858 597454
rect 586302 560898 586858 561454
rect 586302 524898 586858 525454
rect 586302 488898 586858 489454
rect 586302 452898 586858 453454
rect 586302 416898 586858 417454
rect 586302 380898 586858 381454
rect 586302 344898 586858 345454
rect 586302 308898 586858 309454
rect 586302 272898 586858 273454
rect 586302 236898 586858 237454
rect 586302 200898 586858 201454
rect 586302 164898 586858 165454
rect 586302 128898 586858 129454
rect 586302 92898 586858 93454
rect 586302 56898 586858 57454
rect 586302 20898 586858 21454
rect 586302 -1862 586858 -1306
rect 587262 690618 587818 691174
rect 587262 654618 587818 655174
rect 587262 618618 587818 619174
rect 587262 582618 587818 583174
rect 587262 546618 587818 547174
rect 587262 510618 587818 511174
rect 587262 474618 587818 475174
rect 587262 438618 587818 439174
rect 587262 402618 587818 403174
rect 587262 366618 587818 367174
rect 587262 330618 587818 331174
rect 587262 294618 587818 295174
rect 587262 258618 587818 259174
rect 587262 222618 587818 223174
rect 587262 186618 587818 187174
rect 587262 150618 587818 151174
rect 587262 114618 587818 115174
rect 587262 78618 587818 79174
rect 587262 42618 587818 43174
rect 587262 6618 587818 7174
rect 581546 -2822 582102 -2266
rect 587262 -2822 587818 -2266
rect 588222 672618 588778 673174
rect 588222 636618 588778 637174
rect 588222 600618 588778 601174
rect 588222 564618 588778 565174
rect 588222 528618 588778 529174
rect 588222 492618 588778 493174
rect 588222 456618 588778 457174
rect 588222 420618 588778 421174
rect 588222 384618 588778 385174
rect 588222 348618 588778 349174
rect 588222 312618 588778 313174
rect 588222 276618 588778 277174
rect 588222 240618 588778 241174
rect 588222 204618 588778 205174
rect 588222 168618 588778 169174
rect 588222 132618 588778 133174
rect 588222 96618 588778 97174
rect 588222 60618 588778 61174
rect 588222 24618 588778 25174
rect 588222 -3782 588778 -3226
rect 589182 694338 589738 694894
rect 589182 658338 589738 658894
rect 589182 622338 589738 622894
rect 589182 586338 589738 586894
rect 589182 550338 589738 550894
rect 589182 514338 589738 514894
rect 589182 478338 589738 478894
rect 589182 442338 589738 442894
rect 589182 406338 589738 406894
rect 589182 370338 589738 370894
rect 589182 334338 589738 334894
rect 589182 298338 589738 298894
rect 589182 262338 589738 262894
rect 589182 226338 589738 226894
rect 589182 190338 589738 190894
rect 589182 154338 589738 154894
rect 589182 118338 589738 118894
rect 589182 82338 589738 82894
rect 589182 46338 589738 46894
rect 589182 10338 589738 10894
rect 589182 -4742 589738 -4186
rect 590142 676338 590698 676894
rect 590142 640338 590698 640894
rect 590142 604338 590698 604894
rect 590142 568338 590698 568894
rect 590142 532338 590698 532894
rect 590142 496338 590698 496894
rect 590142 460338 590698 460894
rect 590142 424338 590698 424894
rect 590142 388338 590698 388894
rect 590142 352338 590698 352894
rect 590142 316338 590698 316894
rect 590142 280338 590698 280894
rect 590142 244338 590698 244894
rect 590142 208338 590698 208894
rect 590142 172338 590698 172894
rect 590142 136338 590698 136894
rect 590142 100338 590698 100894
rect 590142 64338 590698 64894
rect 590142 28338 590698 28894
rect 590142 -5702 590698 -5146
rect 591102 698058 591658 698614
rect 591102 662058 591658 662614
rect 591102 626058 591658 626614
rect 591102 590058 591658 590614
rect 591102 554058 591658 554614
rect 591102 518058 591658 518614
rect 591102 482058 591658 482614
rect 591102 446058 591658 446614
rect 591102 410058 591658 410614
rect 591102 374058 591658 374614
rect 591102 338058 591658 338614
rect 591102 302058 591658 302614
rect 591102 266058 591658 266614
rect 591102 230058 591658 230614
rect 591102 194058 591658 194614
rect 591102 158058 591658 158614
rect 591102 122058 591658 122614
rect 591102 86058 591658 86614
rect 591102 50058 591658 50614
rect 591102 14058 591658 14614
rect 591102 -6662 591658 -6106
rect 592062 680058 592618 680614
rect 592062 644058 592618 644614
rect 592062 608058 592618 608614
rect 592062 572058 592618 572614
rect 592062 536058 592618 536614
rect 592062 500058 592618 500614
rect 592062 464058 592618 464614
rect 592062 428058 592618 428614
rect 592062 392058 592618 392614
rect 592062 356058 592618 356614
rect 592062 320058 592618 320614
rect 592062 284058 592618 284614
rect 592062 248058 592618 248614
rect 592062 212058 592618 212614
rect 592062 176058 592618 176614
rect 592062 140058 592618 140614
rect 592062 104058 592618 104614
rect 592062 68058 592618 68614
rect 592062 32058 592618 32614
rect 570986 -7622 571542 -7066
rect 592062 -7622 592618 -7066
<< metal5 >>
rect -8726 711558 592650 711590
rect -8726 711002 -8694 711558
rect -8138 711002 30986 711558
rect 31542 711002 66986 711558
rect 67542 711002 102986 711558
rect 103542 711002 138986 711558
rect 139542 711002 174986 711558
rect 175542 711002 210986 711558
rect 211542 711002 246986 711558
rect 247542 711002 282986 711558
rect 283542 711002 318986 711558
rect 319542 711002 354986 711558
rect 355542 711002 390986 711558
rect 391542 711002 426986 711558
rect 427542 711002 462986 711558
rect 463542 711002 498986 711558
rect 499542 711002 534986 711558
rect 535542 711002 570986 711558
rect 571542 711002 592062 711558
rect 592618 711002 592650 711558
rect -8726 710970 592650 711002
rect -7766 710598 591690 710630
rect -7766 710042 -7734 710598
rect -7178 710042 12986 710598
rect 13542 710042 48986 710598
rect 49542 710042 84986 710598
rect 85542 710042 120986 710598
rect 121542 710042 156986 710598
rect 157542 710042 192986 710598
rect 193542 710042 228986 710598
rect 229542 710042 264986 710598
rect 265542 710042 300986 710598
rect 301542 710042 336986 710598
rect 337542 710042 372986 710598
rect 373542 710042 408986 710598
rect 409542 710042 444986 710598
rect 445542 710042 480986 710598
rect 481542 710042 516986 710598
rect 517542 710042 552986 710598
rect 553542 710042 591102 710598
rect 591658 710042 591690 710598
rect -7766 710010 591690 710042
rect -6806 709638 590730 709670
rect -6806 709082 -6774 709638
rect -6218 709082 27266 709638
rect 27822 709082 63266 709638
rect 63822 709082 99266 709638
rect 99822 709082 135266 709638
rect 135822 709082 171266 709638
rect 171822 709082 207266 709638
rect 207822 709082 243266 709638
rect 243822 709082 279266 709638
rect 279822 709082 315266 709638
rect 315822 709082 351266 709638
rect 351822 709082 387266 709638
rect 387822 709082 423266 709638
rect 423822 709082 459266 709638
rect 459822 709082 495266 709638
rect 495822 709082 531266 709638
rect 531822 709082 567266 709638
rect 567822 709082 590142 709638
rect 590698 709082 590730 709638
rect -6806 709050 590730 709082
rect -5846 708678 589770 708710
rect -5846 708122 -5814 708678
rect -5258 708122 9266 708678
rect 9822 708122 45266 708678
rect 45822 708122 81266 708678
rect 81822 708122 117266 708678
rect 117822 708122 153266 708678
rect 153822 708122 189266 708678
rect 189822 708122 225266 708678
rect 225822 708122 261266 708678
rect 261822 708122 297266 708678
rect 297822 708122 333266 708678
rect 333822 708122 369266 708678
rect 369822 708122 405266 708678
rect 405822 708122 441266 708678
rect 441822 708122 477266 708678
rect 477822 708122 513266 708678
rect 513822 708122 549266 708678
rect 549822 708122 589182 708678
rect 589738 708122 589770 708678
rect -5846 708090 589770 708122
rect -4886 707718 588810 707750
rect -4886 707162 -4854 707718
rect -4298 707162 23546 707718
rect 24102 707162 59546 707718
rect 60102 707162 95546 707718
rect 96102 707162 131546 707718
rect 132102 707162 167546 707718
rect 168102 707162 203546 707718
rect 204102 707162 239546 707718
rect 240102 707162 275546 707718
rect 276102 707162 311546 707718
rect 312102 707162 347546 707718
rect 348102 707162 383546 707718
rect 384102 707162 419546 707718
rect 420102 707162 455546 707718
rect 456102 707162 491546 707718
rect 492102 707162 527546 707718
rect 528102 707162 563546 707718
rect 564102 707162 588222 707718
rect 588778 707162 588810 707718
rect -4886 707130 588810 707162
rect -3926 706758 587850 706790
rect -3926 706202 -3894 706758
rect -3338 706202 5546 706758
rect 6102 706202 41546 706758
rect 42102 706202 77546 706758
rect 78102 706202 113546 706758
rect 114102 706202 149546 706758
rect 150102 706202 185546 706758
rect 186102 706202 221546 706758
rect 222102 706202 257546 706758
rect 258102 706202 293546 706758
rect 294102 706202 329546 706758
rect 330102 706202 365546 706758
rect 366102 706202 401546 706758
rect 402102 706202 437546 706758
rect 438102 706202 473546 706758
rect 474102 706202 509546 706758
rect 510102 706202 545546 706758
rect 546102 706202 581546 706758
rect 582102 706202 587262 706758
rect 587818 706202 587850 706758
rect -3926 706170 587850 706202
rect -2966 705798 586890 705830
rect -2966 705242 -2934 705798
rect -2378 705242 19826 705798
rect 20382 705242 55826 705798
rect 56382 705242 91826 705798
rect 92382 705242 127826 705798
rect 128382 705242 163826 705798
rect 164382 705242 199826 705798
rect 200382 705242 235826 705798
rect 236382 705242 271826 705798
rect 272382 705242 307826 705798
rect 308382 705242 343826 705798
rect 344382 705242 379826 705798
rect 380382 705242 415826 705798
rect 416382 705242 451826 705798
rect 452382 705242 487826 705798
rect 488382 705242 523826 705798
rect 524382 705242 559826 705798
rect 560382 705242 586302 705798
rect 586858 705242 586890 705798
rect -2966 705210 586890 705242
rect -2006 704838 585930 704870
rect -2006 704282 -1974 704838
rect -1418 704282 1826 704838
rect 2382 704282 37826 704838
rect 38382 704282 73826 704838
rect 74382 704282 109826 704838
rect 110382 704282 145826 704838
rect 146382 704282 181826 704838
rect 182382 704282 217826 704838
rect 218382 704282 253826 704838
rect 254382 704282 289826 704838
rect 290382 704282 325826 704838
rect 326382 704282 361826 704838
rect 362382 704282 397826 704838
rect 398382 704282 433826 704838
rect 434382 704282 469826 704838
rect 470382 704282 505826 704838
rect 506382 704282 541826 704838
rect 542382 704282 577826 704838
rect 578382 704282 585342 704838
rect 585898 704282 585930 704838
rect -2006 704250 585930 704282
rect -8726 698614 592650 698646
rect -8726 698058 -7734 698614
rect -7178 698058 12986 698614
rect 13542 698058 48986 698614
rect 49542 698058 84986 698614
rect 85542 698058 120986 698614
rect 121542 698058 156986 698614
rect 157542 698058 192986 698614
rect 193542 698058 228986 698614
rect 229542 698058 264986 698614
rect 265542 698058 300986 698614
rect 301542 698058 336986 698614
rect 337542 698058 372986 698614
rect 373542 698058 408986 698614
rect 409542 698058 444986 698614
rect 445542 698058 480986 698614
rect 481542 698058 516986 698614
rect 517542 698058 552986 698614
rect 553542 698058 591102 698614
rect 591658 698058 592650 698614
rect -8726 698026 592650 698058
rect -6806 694894 590730 694926
rect -6806 694338 -5814 694894
rect -5258 694338 9266 694894
rect 9822 694338 45266 694894
rect 45822 694338 81266 694894
rect 81822 694338 117266 694894
rect 117822 694338 153266 694894
rect 153822 694338 189266 694894
rect 189822 694338 225266 694894
rect 225822 694338 261266 694894
rect 261822 694338 297266 694894
rect 297822 694338 333266 694894
rect 333822 694338 369266 694894
rect 369822 694338 405266 694894
rect 405822 694338 441266 694894
rect 441822 694338 477266 694894
rect 477822 694338 513266 694894
rect 513822 694338 549266 694894
rect 549822 694338 589182 694894
rect 589738 694338 590730 694894
rect -6806 694306 590730 694338
rect -4886 691174 588810 691206
rect -4886 690618 -3894 691174
rect -3338 690618 5546 691174
rect 6102 690618 41546 691174
rect 42102 690618 77546 691174
rect 78102 690618 113546 691174
rect 114102 690618 149546 691174
rect 150102 690618 185546 691174
rect 186102 690618 221546 691174
rect 222102 690618 257546 691174
rect 258102 690618 293546 691174
rect 294102 690618 329546 691174
rect 330102 690618 365546 691174
rect 366102 690618 401546 691174
rect 402102 690618 437546 691174
rect 438102 690618 473546 691174
rect 474102 690618 509546 691174
rect 510102 690618 545546 691174
rect 546102 690618 581546 691174
rect 582102 690618 587262 691174
rect 587818 690618 588810 691174
rect -4886 690586 588810 690618
rect -2966 687454 586890 687486
rect -2966 686898 -1974 687454
rect -1418 686898 1826 687454
rect 2382 686898 37826 687454
rect 38382 686898 73826 687454
rect 74382 686898 109826 687454
rect 110382 686898 145826 687454
rect 146382 686898 181826 687454
rect 182382 686898 217826 687454
rect 218382 686898 253826 687454
rect 254382 686898 289826 687454
rect 290382 686898 325826 687454
rect 326382 686898 361826 687454
rect 362382 686898 397826 687454
rect 398382 686898 433826 687454
rect 434382 686898 469826 687454
rect 470382 686898 505826 687454
rect 506382 686898 541826 687454
rect 542382 686898 577826 687454
rect 578382 686898 585342 687454
rect 585898 686898 586890 687454
rect -2966 686866 586890 686898
rect -8726 680614 592650 680646
rect -8726 680058 -8694 680614
rect -8138 680058 30986 680614
rect 31542 680058 66986 680614
rect 67542 680058 102986 680614
rect 103542 680058 138986 680614
rect 139542 680058 174986 680614
rect 175542 680058 210986 680614
rect 211542 680058 246986 680614
rect 247542 680058 282986 680614
rect 283542 680058 318986 680614
rect 319542 680058 354986 680614
rect 355542 680058 390986 680614
rect 391542 680058 426986 680614
rect 427542 680058 462986 680614
rect 463542 680058 498986 680614
rect 499542 680058 534986 680614
rect 535542 680058 570986 680614
rect 571542 680058 592062 680614
rect 592618 680058 592650 680614
rect -8726 680026 592650 680058
rect -6806 676894 590730 676926
rect -6806 676338 -6774 676894
rect -6218 676338 27266 676894
rect 27822 676338 63266 676894
rect 63822 676338 99266 676894
rect 99822 676338 135266 676894
rect 135822 676338 171266 676894
rect 171822 676338 207266 676894
rect 207822 676338 243266 676894
rect 243822 676338 279266 676894
rect 279822 676338 315266 676894
rect 315822 676338 351266 676894
rect 351822 676338 387266 676894
rect 387822 676338 423266 676894
rect 423822 676338 459266 676894
rect 459822 676338 495266 676894
rect 495822 676338 531266 676894
rect 531822 676338 567266 676894
rect 567822 676338 590142 676894
rect 590698 676338 590730 676894
rect -6806 676306 590730 676338
rect -4886 673174 588810 673206
rect -4886 672618 -4854 673174
rect -4298 672618 23546 673174
rect 24102 672618 59546 673174
rect 60102 672618 95546 673174
rect 96102 672618 131546 673174
rect 132102 672618 167546 673174
rect 168102 672618 203546 673174
rect 204102 672618 239546 673174
rect 240102 672618 275546 673174
rect 276102 672618 311546 673174
rect 312102 672618 347546 673174
rect 348102 672618 383546 673174
rect 384102 672618 419546 673174
rect 420102 672618 455546 673174
rect 456102 672618 491546 673174
rect 492102 672618 527546 673174
rect 528102 672618 563546 673174
rect 564102 672618 588222 673174
rect 588778 672618 588810 673174
rect -4886 672586 588810 672618
rect -2966 669454 586890 669486
rect -2966 668898 -2934 669454
rect -2378 668898 19826 669454
rect 20382 668898 55826 669454
rect 56382 668898 91826 669454
rect 92382 668898 127826 669454
rect 128382 668898 163826 669454
rect 164382 668898 199826 669454
rect 200382 668898 235826 669454
rect 236382 668898 271826 669454
rect 272382 668898 307826 669454
rect 308382 668898 343826 669454
rect 344382 668898 379826 669454
rect 380382 668898 415826 669454
rect 416382 668898 451826 669454
rect 452382 668898 487826 669454
rect 488382 668898 523826 669454
rect 524382 668898 559826 669454
rect 560382 668898 586302 669454
rect 586858 668898 586890 669454
rect -2966 668866 586890 668898
rect -8726 662614 592650 662646
rect -8726 662058 -7734 662614
rect -7178 662058 12986 662614
rect 13542 662058 48986 662614
rect 49542 662058 84986 662614
rect 85542 662058 120986 662614
rect 121542 662058 156986 662614
rect 157542 662058 192986 662614
rect 193542 662058 228986 662614
rect 229542 662058 264986 662614
rect 265542 662058 300986 662614
rect 301542 662058 336986 662614
rect 337542 662058 372986 662614
rect 373542 662058 408986 662614
rect 409542 662058 444986 662614
rect 445542 662058 480986 662614
rect 481542 662058 516986 662614
rect 517542 662058 552986 662614
rect 553542 662058 591102 662614
rect 591658 662058 592650 662614
rect -8726 662026 592650 662058
rect -6806 658894 590730 658926
rect -6806 658338 -5814 658894
rect -5258 658338 9266 658894
rect 9822 658338 45266 658894
rect 45822 658338 81266 658894
rect 81822 658338 117266 658894
rect 117822 658338 153266 658894
rect 153822 658338 189266 658894
rect 189822 658338 225266 658894
rect 225822 658338 261266 658894
rect 261822 658338 297266 658894
rect 297822 658338 333266 658894
rect 333822 658338 369266 658894
rect 369822 658338 405266 658894
rect 405822 658338 441266 658894
rect 441822 658338 477266 658894
rect 477822 658338 513266 658894
rect 513822 658338 549266 658894
rect 549822 658338 589182 658894
rect 589738 658338 590730 658894
rect -6806 658306 590730 658338
rect -4886 655174 588810 655206
rect -4886 654618 -3894 655174
rect -3338 654618 5546 655174
rect 6102 654618 41546 655174
rect 42102 654618 77546 655174
rect 78102 654618 113546 655174
rect 114102 654618 149546 655174
rect 150102 654618 185546 655174
rect 186102 654618 221546 655174
rect 222102 654618 257546 655174
rect 258102 654618 293546 655174
rect 294102 654618 329546 655174
rect 330102 654618 365546 655174
rect 366102 654618 401546 655174
rect 402102 654618 437546 655174
rect 438102 654618 473546 655174
rect 474102 654618 509546 655174
rect 510102 654618 545546 655174
rect 546102 654618 581546 655174
rect 582102 654618 587262 655174
rect 587818 654618 588810 655174
rect -4886 654586 588810 654618
rect -2966 651454 586890 651486
rect -2966 650898 -1974 651454
rect -1418 650898 1826 651454
rect 2382 650898 37826 651454
rect 38382 650898 73826 651454
rect 74382 650898 109826 651454
rect 110382 650898 145826 651454
rect 146382 650898 181826 651454
rect 182382 650898 217826 651454
rect 218382 650898 253826 651454
rect 254382 650898 289826 651454
rect 290382 650898 325826 651454
rect 326382 650898 361826 651454
rect 362382 650898 397826 651454
rect 398382 650898 433826 651454
rect 434382 650898 469826 651454
rect 470382 650898 505826 651454
rect 506382 650898 541826 651454
rect 542382 650898 577826 651454
rect 578382 650898 585342 651454
rect 585898 650898 586890 651454
rect -2966 650866 586890 650898
rect -8726 644614 592650 644646
rect -8726 644058 -8694 644614
rect -8138 644058 30986 644614
rect 31542 644058 66986 644614
rect 67542 644058 102986 644614
rect 103542 644058 138986 644614
rect 139542 644058 174986 644614
rect 175542 644058 210986 644614
rect 211542 644058 246986 644614
rect 247542 644058 282986 644614
rect 283542 644058 318986 644614
rect 319542 644058 354986 644614
rect 355542 644058 390986 644614
rect 391542 644058 426986 644614
rect 427542 644058 462986 644614
rect 463542 644058 498986 644614
rect 499542 644058 534986 644614
rect 535542 644058 570986 644614
rect 571542 644058 592062 644614
rect 592618 644058 592650 644614
rect -8726 644026 592650 644058
rect -6806 640894 590730 640926
rect -6806 640338 -6774 640894
rect -6218 640338 27266 640894
rect 27822 640338 63266 640894
rect 63822 640338 99266 640894
rect 99822 640338 135266 640894
rect 135822 640338 171266 640894
rect 171822 640338 207266 640894
rect 207822 640338 243266 640894
rect 243822 640338 279266 640894
rect 279822 640338 315266 640894
rect 315822 640338 351266 640894
rect 351822 640338 387266 640894
rect 387822 640338 423266 640894
rect 423822 640338 459266 640894
rect 459822 640338 495266 640894
rect 495822 640338 531266 640894
rect 531822 640338 567266 640894
rect 567822 640338 590142 640894
rect 590698 640338 590730 640894
rect -6806 640306 590730 640338
rect -4886 637174 588810 637206
rect -4886 636618 -4854 637174
rect -4298 636618 23546 637174
rect 24102 636618 59546 637174
rect 60102 636618 95546 637174
rect 96102 636618 131546 637174
rect 132102 636618 167546 637174
rect 168102 636618 203546 637174
rect 204102 636618 239546 637174
rect 240102 636618 275546 637174
rect 276102 636618 311546 637174
rect 312102 636618 347546 637174
rect 348102 636618 383546 637174
rect 384102 636618 419546 637174
rect 420102 636618 455546 637174
rect 456102 636618 491546 637174
rect 492102 636618 527546 637174
rect 528102 636618 563546 637174
rect 564102 636618 588222 637174
rect 588778 636618 588810 637174
rect -4886 636586 588810 636618
rect -2966 633454 586890 633486
rect -2966 632898 -2934 633454
rect -2378 632898 19826 633454
rect 20382 632898 55826 633454
rect 56382 632898 91826 633454
rect 92382 632898 127826 633454
rect 128382 632898 163826 633454
rect 164382 632898 199826 633454
rect 200382 632898 235826 633454
rect 236382 632898 271826 633454
rect 272382 632898 307826 633454
rect 308382 632898 343826 633454
rect 344382 632898 379826 633454
rect 380382 632898 415826 633454
rect 416382 632898 451826 633454
rect 452382 632898 487826 633454
rect 488382 632898 523826 633454
rect 524382 632898 559826 633454
rect 560382 632898 586302 633454
rect 586858 632898 586890 633454
rect -2966 632866 586890 632898
rect -8726 626614 592650 626646
rect -8726 626058 -7734 626614
rect -7178 626058 12986 626614
rect 13542 626058 48986 626614
rect 49542 626058 84986 626614
rect 85542 626058 120986 626614
rect 121542 626058 156986 626614
rect 157542 626058 192986 626614
rect 193542 626058 228986 626614
rect 229542 626058 264986 626614
rect 265542 626058 300986 626614
rect 301542 626058 336986 626614
rect 337542 626058 372986 626614
rect 373542 626058 408986 626614
rect 409542 626058 444986 626614
rect 445542 626058 480986 626614
rect 481542 626058 516986 626614
rect 517542 626058 552986 626614
rect 553542 626058 591102 626614
rect 591658 626058 592650 626614
rect -8726 626026 592650 626058
rect -6806 622894 590730 622926
rect -6806 622338 -5814 622894
rect -5258 622338 9266 622894
rect 9822 622338 45266 622894
rect 45822 622338 81266 622894
rect 81822 622338 117266 622894
rect 117822 622338 153266 622894
rect 153822 622338 189266 622894
rect 189822 622338 225266 622894
rect 225822 622338 261266 622894
rect 261822 622338 297266 622894
rect 297822 622338 333266 622894
rect 333822 622338 369266 622894
rect 369822 622338 405266 622894
rect 405822 622338 441266 622894
rect 441822 622338 477266 622894
rect 477822 622338 513266 622894
rect 513822 622338 549266 622894
rect 549822 622338 589182 622894
rect 589738 622338 590730 622894
rect -6806 622306 590730 622338
rect -4886 619174 588810 619206
rect -4886 618618 -3894 619174
rect -3338 618618 5546 619174
rect 6102 618618 41546 619174
rect 42102 618618 77546 619174
rect 78102 618618 113546 619174
rect 114102 618618 149546 619174
rect 150102 618618 185546 619174
rect 186102 618618 221546 619174
rect 222102 618618 257546 619174
rect 258102 618618 293546 619174
rect 294102 618618 329546 619174
rect 330102 618618 365546 619174
rect 366102 618618 401546 619174
rect 402102 618618 437546 619174
rect 438102 618618 473546 619174
rect 474102 618618 509546 619174
rect 510102 618618 545546 619174
rect 546102 618618 581546 619174
rect 582102 618618 587262 619174
rect 587818 618618 588810 619174
rect -4886 618586 588810 618618
rect -2966 615454 586890 615486
rect -2966 614898 -1974 615454
rect -1418 614898 1826 615454
rect 2382 614898 37826 615454
rect 38382 614898 73826 615454
rect 74382 614898 109826 615454
rect 110382 614898 145826 615454
rect 146382 614898 181826 615454
rect 182382 614898 217826 615454
rect 218382 614898 253826 615454
rect 254382 614898 289826 615454
rect 290382 614898 325826 615454
rect 326382 614898 361826 615454
rect 362382 614898 397826 615454
rect 398382 614898 433826 615454
rect 434382 614898 469826 615454
rect 470382 614898 505826 615454
rect 506382 614898 541826 615454
rect 542382 614898 577826 615454
rect 578382 614898 585342 615454
rect 585898 614898 586890 615454
rect -2966 614866 586890 614898
rect -8726 608614 592650 608646
rect -8726 608058 -8694 608614
rect -8138 608058 30986 608614
rect 31542 608058 66986 608614
rect 67542 608058 102986 608614
rect 103542 608058 138986 608614
rect 139542 608058 174986 608614
rect 175542 608058 210986 608614
rect 211542 608058 246986 608614
rect 247542 608058 282986 608614
rect 283542 608058 318986 608614
rect 319542 608058 354986 608614
rect 355542 608058 390986 608614
rect 391542 608058 426986 608614
rect 427542 608058 462986 608614
rect 463542 608058 498986 608614
rect 499542 608058 534986 608614
rect 535542 608058 570986 608614
rect 571542 608058 592062 608614
rect 592618 608058 592650 608614
rect -8726 608026 592650 608058
rect -6806 604894 590730 604926
rect -6806 604338 -6774 604894
rect -6218 604338 27266 604894
rect 27822 604338 63266 604894
rect 63822 604338 99266 604894
rect 99822 604338 135266 604894
rect 135822 604338 171266 604894
rect 171822 604338 207266 604894
rect 207822 604338 243266 604894
rect 243822 604338 279266 604894
rect 279822 604338 315266 604894
rect 315822 604338 351266 604894
rect 351822 604338 387266 604894
rect 387822 604338 423266 604894
rect 423822 604338 459266 604894
rect 459822 604338 495266 604894
rect 495822 604338 531266 604894
rect 531822 604338 567266 604894
rect 567822 604338 590142 604894
rect 590698 604338 590730 604894
rect -6806 604306 590730 604338
rect -4886 601174 588810 601206
rect -4886 600618 -4854 601174
rect -4298 600618 23546 601174
rect 24102 600618 59546 601174
rect 60102 600618 95546 601174
rect 96102 600618 131546 601174
rect 132102 600618 167546 601174
rect 168102 600618 203546 601174
rect 204102 600618 239546 601174
rect 240102 600618 275546 601174
rect 276102 600618 311546 601174
rect 312102 600618 347546 601174
rect 348102 600618 383546 601174
rect 384102 600618 419546 601174
rect 420102 600618 455546 601174
rect 456102 600618 491546 601174
rect 492102 600618 527546 601174
rect 528102 600618 563546 601174
rect 564102 600618 588222 601174
rect 588778 600618 588810 601174
rect -4886 600586 588810 600618
rect -2966 597454 586890 597486
rect -2966 596898 -2934 597454
rect -2378 596898 19826 597454
rect 20382 596898 55826 597454
rect 56382 596898 91826 597454
rect 92382 596898 127826 597454
rect 128382 596898 163826 597454
rect 164382 596898 199826 597454
rect 200382 596898 235826 597454
rect 236382 596898 271826 597454
rect 272382 596898 307826 597454
rect 308382 596898 343826 597454
rect 344382 596898 379826 597454
rect 380382 596898 415826 597454
rect 416382 596898 451826 597454
rect 452382 596898 487826 597454
rect 488382 596898 523826 597454
rect 524382 596898 559826 597454
rect 560382 596898 586302 597454
rect 586858 596898 586890 597454
rect -2966 596866 586890 596898
rect -8726 590614 592650 590646
rect -8726 590058 -7734 590614
rect -7178 590058 12986 590614
rect 13542 590058 48986 590614
rect 49542 590058 84986 590614
rect 85542 590058 120986 590614
rect 121542 590058 156986 590614
rect 157542 590058 192986 590614
rect 193542 590058 228986 590614
rect 229542 590058 264986 590614
rect 265542 590058 300986 590614
rect 301542 590058 336986 590614
rect 337542 590058 372986 590614
rect 373542 590058 408986 590614
rect 409542 590058 444986 590614
rect 445542 590058 480986 590614
rect 481542 590058 516986 590614
rect 517542 590058 552986 590614
rect 553542 590058 591102 590614
rect 591658 590058 592650 590614
rect -8726 590026 592650 590058
rect -6806 586894 590730 586926
rect -6806 586338 -5814 586894
rect -5258 586338 9266 586894
rect 9822 586338 45266 586894
rect 45822 586338 81266 586894
rect 81822 586338 117266 586894
rect 117822 586338 153266 586894
rect 153822 586338 189266 586894
rect 189822 586338 225266 586894
rect 225822 586338 261266 586894
rect 261822 586338 297266 586894
rect 297822 586338 333266 586894
rect 333822 586338 369266 586894
rect 369822 586338 405266 586894
rect 405822 586338 441266 586894
rect 441822 586338 477266 586894
rect 477822 586338 513266 586894
rect 513822 586338 549266 586894
rect 549822 586338 589182 586894
rect 589738 586338 590730 586894
rect -6806 586306 590730 586338
rect -4886 583174 588810 583206
rect -4886 582618 -3894 583174
rect -3338 582618 5546 583174
rect 6102 582618 41546 583174
rect 42102 582618 77546 583174
rect 78102 582618 113546 583174
rect 114102 582618 149546 583174
rect 150102 582618 185546 583174
rect 186102 582618 221546 583174
rect 222102 582618 257546 583174
rect 258102 582618 293546 583174
rect 294102 582618 329546 583174
rect 330102 582618 365546 583174
rect 366102 582618 401546 583174
rect 402102 582618 437546 583174
rect 438102 582618 473546 583174
rect 474102 582618 509546 583174
rect 510102 582618 545546 583174
rect 546102 582618 581546 583174
rect 582102 582618 587262 583174
rect 587818 582618 588810 583174
rect -4886 582586 588810 582618
rect -2966 579454 586890 579486
rect -2966 578898 -1974 579454
rect -1418 578898 1826 579454
rect 2382 578898 37826 579454
rect 38382 578898 73826 579454
rect 74382 578898 109826 579454
rect 110382 578898 145826 579454
rect 146382 578898 181826 579454
rect 182382 578898 217826 579454
rect 218382 578898 253826 579454
rect 254382 578898 289826 579454
rect 290382 578898 325826 579454
rect 326382 578898 361826 579454
rect 362382 578898 397826 579454
rect 398382 578898 433826 579454
rect 434382 578898 469826 579454
rect 470382 578898 505826 579454
rect 506382 578898 541826 579454
rect 542382 578898 577826 579454
rect 578382 578898 585342 579454
rect 585898 578898 586890 579454
rect -2966 578866 586890 578898
rect -8726 572614 592650 572646
rect -8726 572058 -8694 572614
rect -8138 572058 30986 572614
rect 31542 572058 66986 572614
rect 67542 572058 102986 572614
rect 103542 572058 138986 572614
rect 139542 572058 174986 572614
rect 175542 572058 210986 572614
rect 211542 572058 246986 572614
rect 247542 572058 282986 572614
rect 283542 572058 318986 572614
rect 319542 572058 354986 572614
rect 355542 572058 390986 572614
rect 391542 572058 426986 572614
rect 427542 572058 462986 572614
rect 463542 572058 498986 572614
rect 499542 572058 534986 572614
rect 535542 572058 570986 572614
rect 571542 572058 592062 572614
rect 592618 572058 592650 572614
rect -8726 572026 592650 572058
rect -6806 568894 590730 568926
rect -6806 568338 -6774 568894
rect -6218 568338 27266 568894
rect 27822 568338 63266 568894
rect 63822 568338 99266 568894
rect 99822 568338 135266 568894
rect 135822 568338 171266 568894
rect 171822 568338 207266 568894
rect 207822 568338 243266 568894
rect 243822 568338 279266 568894
rect 279822 568338 315266 568894
rect 315822 568338 351266 568894
rect 351822 568338 387266 568894
rect 387822 568338 423266 568894
rect 423822 568338 459266 568894
rect 459822 568338 495266 568894
rect 495822 568338 531266 568894
rect 531822 568338 567266 568894
rect 567822 568338 590142 568894
rect 590698 568338 590730 568894
rect -6806 568306 590730 568338
rect -4886 565174 588810 565206
rect -4886 564618 -4854 565174
rect -4298 564618 23546 565174
rect 24102 564618 59546 565174
rect 60102 564618 95546 565174
rect 96102 564618 131546 565174
rect 132102 564618 167546 565174
rect 168102 564618 203546 565174
rect 204102 564618 239546 565174
rect 240102 564618 275546 565174
rect 276102 564618 311546 565174
rect 312102 564618 347546 565174
rect 348102 564618 383546 565174
rect 384102 564618 419546 565174
rect 420102 564618 455546 565174
rect 456102 564618 491546 565174
rect 492102 564618 527546 565174
rect 528102 564618 563546 565174
rect 564102 564618 588222 565174
rect 588778 564618 588810 565174
rect -4886 564586 588810 564618
rect -2966 561454 586890 561486
rect -2966 560898 -2934 561454
rect -2378 560898 19826 561454
rect 20382 560898 55826 561454
rect 56382 560898 91826 561454
rect 92382 560898 127826 561454
rect 128382 560898 163826 561454
rect 164382 560898 199826 561454
rect 200382 560898 235826 561454
rect 236382 560898 271826 561454
rect 272382 560898 307826 561454
rect 308382 560898 343826 561454
rect 344382 560898 379826 561454
rect 380382 560898 415826 561454
rect 416382 560898 451826 561454
rect 452382 560898 487826 561454
rect 488382 560898 523826 561454
rect 524382 560898 559826 561454
rect 560382 560898 586302 561454
rect 586858 560898 586890 561454
rect -2966 560866 586890 560898
rect -8726 554614 592650 554646
rect -8726 554058 -7734 554614
rect -7178 554058 12986 554614
rect 13542 554058 48986 554614
rect 49542 554058 84986 554614
rect 85542 554058 120986 554614
rect 121542 554058 156986 554614
rect 157542 554058 192986 554614
rect 193542 554058 228986 554614
rect 229542 554058 264986 554614
rect 265542 554058 300986 554614
rect 301542 554058 336986 554614
rect 337542 554058 372986 554614
rect 373542 554058 408986 554614
rect 409542 554058 444986 554614
rect 445542 554058 480986 554614
rect 481542 554058 516986 554614
rect 517542 554058 552986 554614
rect 553542 554058 591102 554614
rect 591658 554058 592650 554614
rect -8726 554026 592650 554058
rect -6806 550894 590730 550926
rect -6806 550338 -5814 550894
rect -5258 550338 9266 550894
rect 9822 550338 45266 550894
rect 45822 550338 81266 550894
rect 81822 550338 117266 550894
rect 117822 550338 153266 550894
rect 153822 550338 189266 550894
rect 189822 550338 225266 550894
rect 225822 550338 261266 550894
rect 261822 550338 297266 550894
rect 297822 550338 333266 550894
rect 333822 550338 369266 550894
rect 369822 550338 405266 550894
rect 405822 550338 441266 550894
rect 441822 550338 477266 550894
rect 477822 550338 513266 550894
rect 513822 550338 549266 550894
rect 549822 550338 589182 550894
rect 589738 550338 590730 550894
rect -6806 550306 590730 550338
rect -4886 547174 588810 547206
rect -4886 546618 -3894 547174
rect -3338 546618 5546 547174
rect 6102 546618 41546 547174
rect 42102 546618 77546 547174
rect 78102 546618 113546 547174
rect 114102 546618 149546 547174
rect 150102 546618 185546 547174
rect 186102 546618 221546 547174
rect 222102 546618 257546 547174
rect 258102 546618 293546 547174
rect 294102 546618 329546 547174
rect 330102 546618 365546 547174
rect 366102 546618 401546 547174
rect 402102 546618 437546 547174
rect 438102 546618 473546 547174
rect 474102 546618 509546 547174
rect 510102 546618 545546 547174
rect 546102 546618 581546 547174
rect 582102 546618 587262 547174
rect 587818 546618 588810 547174
rect -4886 546586 588810 546618
rect -2966 543454 586890 543486
rect -2966 542898 -1974 543454
rect -1418 542898 1826 543454
rect 2382 542898 37826 543454
rect 38382 542898 73826 543454
rect 74382 542898 109826 543454
rect 110382 542898 145826 543454
rect 146382 542898 181826 543454
rect 182382 542898 217826 543454
rect 218382 542898 253826 543454
rect 254382 542898 289826 543454
rect 290382 542898 325826 543454
rect 326382 542898 361826 543454
rect 362382 542898 397826 543454
rect 398382 542898 433826 543454
rect 434382 542898 469826 543454
rect 470382 542898 505826 543454
rect 506382 542898 541826 543454
rect 542382 542898 577826 543454
rect 578382 542898 585342 543454
rect 585898 542898 586890 543454
rect -2966 542866 586890 542898
rect -8726 536614 592650 536646
rect -8726 536058 -8694 536614
rect -8138 536058 30986 536614
rect 31542 536058 66986 536614
rect 67542 536058 102986 536614
rect 103542 536058 138986 536614
rect 139542 536058 174986 536614
rect 175542 536058 210986 536614
rect 211542 536058 246986 536614
rect 247542 536058 282986 536614
rect 283542 536058 318986 536614
rect 319542 536058 354986 536614
rect 355542 536058 390986 536614
rect 391542 536058 426986 536614
rect 427542 536058 462986 536614
rect 463542 536058 498986 536614
rect 499542 536058 534986 536614
rect 535542 536058 570986 536614
rect 571542 536058 592062 536614
rect 592618 536058 592650 536614
rect -8726 536026 592650 536058
rect -6806 532894 590730 532926
rect -6806 532338 -6774 532894
rect -6218 532338 27266 532894
rect 27822 532338 63266 532894
rect 63822 532338 99266 532894
rect 99822 532338 135266 532894
rect 135822 532338 171266 532894
rect 171822 532338 207266 532894
rect 207822 532338 243266 532894
rect 243822 532338 279266 532894
rect 279822 532338 315266 532894
rect 315822 532338 351266 532894
rect 351822 532338 387266 532894
rect 387822 532338 423266 532894
rect 423822 532338 459266 532894
rect 459822 532338 495266 532894
rect 495822 532338 531266 532894
rect 531822 532338 567266 532894
rect 567822 532338 590142 532894
rect 590698 532338 590730 532894
rect -6806 532306 590730 532338
rect -4886 529174 588810 529206
rect -4886 528618 -4854 529174
rect -4298 528618 23546 529174
rect 24102 528618 59546 529174
rect 60102 528618 95546 529174
rect 96102 528618 131546 529174
rect 132102 528618 167546 529174
rect 168102 528618 203546 529174
rect 204102 528618 239546 529174
rect 240102 528618 275546 529174
rect 276102 528618 311546 529174
rect 312102 528618 347546 529174
rect 348102 528618 383546 529174
rect 384102 528618 419546 529174
rect 420102 528618 455546 529174
rect 456102 528618 491546 529174
rect 492102 528618 527546 529174
rect 528102 528618 563546 529174
rect 564102 528618 588222 529174
rect 588778 528618 588810 529174
rect -4886 528586 588810 528618
rect -2966 525454 586890 525486
rect -2966 524898 -2934 525454
rect -2378 524898 19826 525454
rect 20382 524898 55826 525454
rect 56382 524898 91826 525454
rect 92382 524898 127826 525454
rect 128382 524898 163826 525454
rect 164382 524898 199826 525454
rect 200382 524898 235826 525454
rect 236382 524898 271826 525454
rect 272382 524898 307826 525454
rect 308382 524898 343826 525454
rect 344382 524898 379826 525454
rect 380382 524898 415826 525454
rect 416382 524898 451826 525454
rect 452382 524898 487826 525454
rect 488382 524898 523826 525454
rect 524382 524898 559826 525454
rect 560382 524898 586302 525454
rect 586858 524898 586890 525454
rect -2966 524866 586890 524898
rect -8726 518614 592650 518646
rect -8726 518058 -7734 518614
rect -7178 518058 12986 518614
rect 13542 518058 48986 518614
rect 49542 518058 84986 518614
rect 85542 518058 120986 518614
rect 121542 518058 156986 518614
rect 157542 518058 192986 518614
rect 193542 518058 228986 518614
rect 229542 518058 264986 518614
rect 265542 518058 300986 518614
rect 301542 518058 336986 518614
rect 337542 518058 372986 518614
rect 373542 518058 408986 518614
rect 409542 518058 444986 518614
rect 445542 518058 480986 518614
rect 481542 518058 516986 518614
rect 517542 518058 552986 518614
rect 553542 518058 591102 518614
rect 591658 518058 592650 518614
rect -8726 518026 592650 518058
rect -6806 514894 590730 514926
rect -6806 514338 -5814 514894
rect -5258 514338 9266 514894
rect 9822 514338 45266 514894
rect 45822 514338 81266 514894
rect 81822 514338 117266 514894
rect 117822 514338 153266 514894
rect 153822 514338 189266 514894
rect 189822 514338 225266 514894
rect 225822 514338 261266 514894
rect 261822 514338 297266 514894
rect 297822 514338 333266 514894
rect 333822 514338 369266 514894
rect 369822 514338 405266 514894
rect 405822 514338 441266 514894
rect 441822 514338 477266 514894
rect 477822 514338 513266 514894
rect 513822 514338 549266 514894
rect 549822 514338 589182 514894
rect 589738 514338 590730 514894
rect -6806 514306 590730 514338
rect -4886 511174 588810 511206
rect -4886 510618 -3894 511174
rect -3338 510618 5546 511174
rect 6102 510618 41546 511174
rect 42102 510618 77546 511174
rect 78102 510618 113546 511174
rect 114102 510618 149546 511174
rect 150102 510618 185546 511174
rect 186102 510618 221546 511174
rect 222102 510618 257546 511174
rect 258102 510618 293546 511174
rect 294102 510618 329546 511174
rect 330102 510618 365546 511174
rect 366102 510618 401546 511174
rect 402102 510618 437546 511174
rect 438102 510618 473546 511174
rect 474102 510618 509546 511174
rect 510102 510618 545546 511174
rect 546102 510618 581546 511174
rect 582102 510618 587262 511174
rect 587818 510618 588810 511174
rect -4886 510586 588810 510618
rect -2966 507454 586890 507486
rect -2966 506898 -1974 507454
rect -1418 506898 1826 507454
rect 2382 506898 37826 507454
rect 38382 506898 73826 507454
rect 74382 506898 109826 507454
rect 110382 506898 145826 507454
rect 146382 506898 181826 507454
rect 182382 506898 217826 507454
rect 218382 506898 253826 507454
rect 254382 506898 289826 507454
rect 290382 506898 325826 507454
rect 326382 506898 361826 507454
rect 362382 506898 397826 507454
rect 398382 506898 433826 507454
rect 434382 506898 469826 507454
rect 470382 506898 505826 507454
rect 506382 506898 541826 507454
rect 542382 506898 577826 507454
rect 578382 506898 585342 507454
rect 585898 506898 586890 507454
rect -2966 506866 586890 506898
rect -8726 500614 592650 500646
rect -8726 500058 -8694 500614
rect -8138 500058 30986 500614
rect 31542 500058 66986 500614
rect 67542 500058 102986 500614
rect 103542 500058 138986 500614
rect 139542 500058 174986 500614
rect 175542 500058 210986 500614
rect 211542 500058 246986 500614
rect 247542 500058 282986 500614
rect 283542 500058 318986 500614
rect 319542 500058 354986 500614
rect 355542 500058 390986 500614
rect 391542 500058 426986 500614
rect 427542 500058 462986 500614
rect 463542 500058 498986 500614
rect 499542 500058 534986 500614
rect 535542 500058 570986 500614
rect 571542 500058 592062 500614
rect 592618 500058 592650 500614
rect -8726 500026 592650 500058
rect -6806 496894 590730 496926
rect -6806 496338 -6774 496894
rect -6218 496338 27266 496894
rect 27822 496338 63266 496894
rect 63822 496338 99266 496894
rect 99822 496338 135266 496894
rect 135822 496338 171266 496894
rect 171822 496338 207266 496894
rect 207822 496338 243266 496894
rect 243822 496338 279266 496894
rect 279822 496338 315266 496894
rect 315822 496338 351266 496894
rect 351822 496338 387266 496894
rect 387822 496338 423266 496894
rect 423822 496338 459266 496894
rect 459822 496338 495266 496894
rect 495822 496338 531266 496894
rect 531822 496338 567266 496894
rect 567822 496338 590142 496894
rect 590698 496338 590730 496894
rect -6806 496306 590730 496338
rect -4886 493174 588810 493206
rect -4886 492618 -4854 493174
rect -4298 492618 23546 493174
rect 24102 492618 59546 493174
rect 60102 492618 95546 493174
rect 96102 492618 131546 493174
rect 132102 492618 167546 493174
rect 168102 492618 203546 493174
rect 204102 492618 239546 493174
rect 240102 492618 275546 493174
rect 276102 492618 311546 493174
rect 312102 492618 347546 493174
rect 348102 492618 383546 493174
rect 384102 492618 419546 493174
rect 420102 492618 455546 493174
rect 456102 492618 491546 493174
rect 492102 492618 527546 493174
rect 528102 492618 563546 493174
rect 564102 492618 588222 493174
rect 588778 492618 588810 493174
rect -4886 492586 588810 492618
rect -2966 489454 586890 489486
rect -2966 488898 -2934 489454
rect -2378 488898 19826 489454
rect 20382 488898 55826 489454
rect 56382 488898 91826 489454
rect 92382 488898 127826 489454
rect 128382 488898 163826 489454
rect 164382 488898 199826 489454
rect 200382 488898 415826 489454
rect 416382 488898 451826 489454
rect 452382 488898 487826 489454
rect 488382 488898 523826 489454
rect 524382 488898 559826 489454
rect 560382 488898 586302 489454
rect 586858 488898 586890 489454
rect -2966 488866 586890 488898
rect -8726 482614 592650 482646
rect -8726 482058 -7734 482614
rect -7178 482058 12986 482614
rect 13542 482058 48986 482614
rect 49542 482058 84986 482614
rect 85542 482058 120986 482614
rect 121542 482058 156986 482614
rect 157542 482058 192986 482614
rect 193542 482058 228986 482614
rect 229542 482058 408986 482614
rect 409542 482058 444986 482614
rect 445542 482058 480986 482614
rect 481542 482058 516986 482614
rect 517542 482058 552986 482614
rect 553542 482058 591102 482614
rect 591658 482058 592650 482614
rect -8726 482026 592650 482058
rect -6806 478894 590730 478926
rect -6806 478338 -5814 478894
rect -5258 478338 9266 478894
rect 9822 478338 45266 478894
rect 45822 478338 81266 478894
rect 81822 478338 117266 478894
rect 117822 478338 153266 478894
rect 153822 478338 189266 478894
rect 189822 478338 225266 478894
rect 225822 478338 405266 478894
rect 405822 478338 441266 478894
rect 441822 478338 477266 478894
rect 477822 478338 513266 478894
rect 513822 478338 549266 478894
rect 549822 478338 589182 478894
rect 589738 478338 590730 478894
rect -6806 478306 590730 478338
rect -4886 475174 588810 475206
rect -4886 474618 -3894 475174
rect -3338 474618 5546 475174
rect 6102 474618 41546 475174
rect 42102 474618 77546 475174
rect 78102 474618 113546 475174
rect 114102 474618 149546 475174
rect 150102 474618 185546 475174
rect 186102 474618 221546 475174
rect 222102 474618 401546 475174
rect 402102 474618 437546 475174
rect 438102 474618 473546 475174
rect 474102 474618 509546 475174
rect 510102 474618 545546 475174
rect 546102 474618 581546 475174
rect 582102 474618 587262 475174
rect 587818 474618 588810 475174
rect -4886 474586 588810 474618
rect -2966 471454 586890 471486
rect -2966 470898 -1974 471454
rect -1418 470898 1826 471454
rect 2382 470898 37826 471454
rect 38382 470898 73826 471454
rect 74382 470898 109826 471454
rect 110382 470898 145826 471454
rect 146382 470898 181826 471454
rect 182382 470898 217826 471454
rect 218382 471218 239250 471454
rect 239486 471218 269970 471454
rect 270206 471218 300690 471454
rect 300926 471218 331410 471454
rect 331646 471218 362130 471454
rect 362366 471218 397826 471454
rect 218382 471134 397826 471218
rect 218382 470898 239250 471134
rect 239486 470898 269970 471134
rect 270206 470898 300690 471134
rect 300926 470898 331410 471134
rect 331646 470898 362130 471134
rect 362366 470898 397826 471134
rect 398382 470898 433826 471454
rect 434382 470898 469826 471454
rect 470382 470898 505826 471454
rect 506382 470898 541826 471454
rect 542382 470898 577826 471454
rect 578382 470898 585342 471454
rect 585898 470898 586890 471454
rect -2966 470866 586890 470898
rect -8726 464614 592650 464646
rect -8726 464058 -8694 464614
rect -8138 464058 30986 464614
rect 31542 464058 66986 464614
rect 67542 464058 102986 464614
rect 103542 464058 138986 464614
rect 139542 464058 174986 464614
rect 175542 464058 210986 464614
rect 211542 464058 390986 464614
rect 391542 464058 426986 464614
rect 427542 464058 462986 464614
rect 463542 464058 498986 464614
rect 499542 464058 534986 464614
rect 535542 464058 570986 464614
rect 571542 464058 592062 464614
rect 592618 464058 592650 464614
rect -8726 464026 592650 464058
rect -6806 460894 590730 460926
rect -6806 460338 -6774 460894
rect -6218 460338 27266 460894
rect 27822 460338 63266 460894
rect 63822 460338 99266 460894
rect 99822 460338 135266 460894
rect 135822 460338 171266 460894
rect 171822 460338 207266 460894
rect 207822 460338 387266 460894
rect 387822 460338 423266 460894
rect 423822 460338 459266 460894
rect 459822 460338 495266 460894
rect 495822 460338 531266 460894
rect 531822 460338 567266 460894
rect 567822 460338 590142 460894
rect 590698 460338 590730 460894
rect -6806 460306 590730 460338
rect -4886 457174 588810 457206
rect -4886 456618 -4854 457174
rect -4298 456618 23546 457174
rect 24102 456618 59546 457174
rect 60102 456618 95546 457174
rect 96102 456618 131546 457174
rect 132102 456618 167546 457174
rect 168102 456618 203546 457174
rect 204102 456618 419546 457174
rect 420102 456618 455546 457174
rect 456102 456618 491546 457174
rect 492102 456618 527546 457174
rect 528102 456618 563546 457174
rect 564102 456618 588222 457174
rect 588778 456618 588810 457174
rect -4886 456586 588810 456618
rect -2966 453454 586890 453486
rect -2966 452898 -2934 453454
rect -2378 452898 19826 453454
rect 20382 452898 55826 453454
rect 56382 452898 91826 453454
rect 92382 452898 127826 453454
rect 128382 452898 163826 453454
rect 164382 452898 199826 453454
rect 200382 453218 254610 453454
rect 254846 453218 285330 453454
rect 285566 453218 316050 453454
rect 316286 453218 346770 453454
rect 347006 453218 377490 453454
rect 377726 453218 415826 453454
rect 200382 453134 415826 453218
rect 200382 452898 254610 453134
rect 254846 452898 285330 453134
rect 285566 452898 316050 453134
rect 316286 452898 346770 453134
rect 347006 452898 377490 453134
rect 377726 452898 415826 453134
rect 416382 452898 451826 453454
rect 452382 452898 487826 453454
rect 488382 452898 523826 453454
rect 524382 452898 559826 453454
rect 560382 452898 586302 453454
rect 586858 452898 586890 453454
rect -2966 452866 586890 452898
rect -8726 446614 592650 446646
rect -8726 446058 -7734 446614
rect -7178 446058 12986 446614
rect 13542 446058 48986 446614
rect 49542 446058 84986 446614
rect 85542 446058 120986 446614
rect 121542 446058 156986 446614
rect 157542 446058 192986 446614
rect 193542 446058 228986 446614
rect 229542 446058 408986 446614
rect 409542 446058 444986 446614
rect 445542 446058 480986 446614
rect 481542 446058 516986 446614
rect 517542 446058 552986 446614
rect 553542 446058 591102 446614
rect 591658 446058 592650 446614
rect -8726 446026 592650 446058
rect -6806 442894 590730 442926
rect -6806 442338 -5814 442894
rect -5258 442338 9266 442894
rect 9822 442338 45266 442894
rect 45822 442338 81266 442894
rect 81822 442338 117266 442894
rect 117822 442338 153266 442894
rect 153822 442338 189266 442894
rect 189822 442338 225266 442894
rect 225822 442338 405266 442894
rect 405822 442338 441266 442894
rect 441822 442338 477266 442894
rect 477822 442338 513266 442894
rect 513822 442338 549266 442894
rect 549822 442338 589182 442894
rect 589738 442338 590730 442894
rect -6806 442306 590730 442338
rect -4886 439174 588810 439206
rect -4886 438618 -3894 439174
rect -3338 438618 5546 439174
rect 6102 438618 41546 439174
rect 42102 438618 77546 439174
rect 78102 438618 113546 439174
rect 114102 438618 149546 439174
rect 150102 438618 185546 439174
rect 186102 438618 221546 439174
rect 222102 438618 401546 439174
rect 402102 438618 437546 439174
rect 438102 438618 473546 439174
rect 474102 438618 509546 439174
rect 510102 438618 545546 439174
rect 546102 438618 581546 439174
rect 582102 438618 587262 439174
rect 587818 438618 588810 439174
rect -4886 438586 588810 438618
rect -2966 435454 586890 435486
rect -2966 434898 -1974 435454
rect -1418 434898 1826 435454
rect 2382 434898 37826 435454
rect 38382 434898 73826 435454
rect 74382 434898 109826 435454
rect 110382 434898 145826 435454
rect 146382 434898 181826 435454
rect 182382 434898 217826 435454
rect 218382 435218 239250 435454
rect 239486 435218 269970 435454
rect 270206 435218 300690 435454
rect 300926 435218 331410 435454
rect 331646 435218 362130 435454
rect 362366 435218 397826 435454
rect 218382 435134 397826 435218
rect 218382 434898 239250 435134
rect 239486 434898 269970 435134
rect 270206 434898 300690 435134
rect 300926 434898 331410 435134
rect 331646 434898 362130 435134
rect 362366 434898 397826 435134
rect 398382 434898 433826 435454
rect 434382 434898 469826 435454
rect 470382 434898 505826 435454
rect 506382 434898 541826 435454
rect 542382 434898 577826 435454
rect 578382 434898 585342 435454
rect 585898 434898 586890 435454
rect -2966 434866 586890 434898
rect -8726 428614 592650 428646
rect -8726 428058 -8694 428614
rect -8138 428058 30986 428614
rect 31542 428058 66986 428614
rect 67542 428058 102986 428614
rect 103542 428058 138986 428614
rect 139542 428058 174986 428614
rect 175542 428058 210986 428614
rect 211542 428058 390986 428614
rect 391542 428058 426986 428614
rect 427542 428058 462986 428614
rect 463542 428058 498986 428614
rect 499542 428058 534986 428614
rect 535542 428058 570986 428614
rect 571542 428058 592062 428614
rect 592618 428058 592650 428614
rect -8726 428026 592650 428058
rect -6806 424894 590730 424926
rect -6806 424338 -6774 424894
rect -6218 424338 27266 424894
rect 27822 424338 63266 424894
rect 63822 424338 99266 424894
rect 99822 424338 135266 424894
rect 135822 424338 171266 424894
rect 171822 424338 207266 424894
rect 207822 424338 387266 424894
rect 387822 424338 423266 424894
rect 423822 424338 459266 424894
rect 459822 424338 495266 424894
rect 495822 424338 531266 424894
rect 531822 424338 567266 424894
rect 567822 424338 590142 424894
rect 590698 424338 590730 424894
rect -6806 424306 590730 424338
rect -4886 421174 588810 421206
rect -4886 420618 -4854 421174
rect -4298 420618 23546 421174
rect 24102 420618 59546 421174
rect 60102 420618 95546 421174
rect 96102 420618 131546 421174
rect 132102 420618 167546 421174
rect 168102 420618 203546 421174
rect 204102 420618 419546 421174
rect 420102 420618 455546 421174
rect 456102 420618 491546 421174
rect 492102 420618 527546 421174
rect 528102 420618 563546 421174
rect 564102 420618 588222 421174
rect 588778 420618 588810 421174
rect -4886 420586 588810 420618
rect -2966 417454 586890 417486
rect -2966 416898 -2934 417454
rect -2378 416898 19826 417454
rect 20382 416898 55826 417454
rect 56382 416898 91826 417454
rect 92382 416898 127826 417454
rect 128382 416898 163826 417454
rect 164382 416898 199826 417454
rect 200382 417218 254610 417454
rect 254846 417218 285330 417454
rect 285566 417218 316050 417454
rect 316286 417218 346770 417454
rect 347006 417218 377490 417454
rect 377726 417218 415826 417454
rect 200382 417134 415826 417218
rect 200382 416898 254610 417134
rect 254846 416898 285330 417134
rect 285566 416898 316050 417134
rect 316286 416898 346770 417134
rect 347006 416898 377490 417134
rect 377726 416898 415826 417134
rect 416382 416898 451826 417454
rect 452382 416898 487826 417454
rect 488382 416898 523826 417454
rect 524382 416898 559826 417454
rect 560382 416898 586302 417454
rect 586858 416898 586890 417454
rect -2966 416866 586890 416898
rect -8726 410614 592650 410646
rect -8726 410058 -7734 410614
rect -7178 410058 12986 410614
rect 13542 410058 48986 410614
rect 49542 410058 84986 410614
rect 85542 410058 120986 410614
rect 121542 410058 156986 410614
rect 157542 410058 192986 410614
rect 193542 410058 228986 410614
rect 229542 410058 408986 410614
rect 409542 410058 444986 410614
rect 445542 410058 480986 410614
rect 481542 410058 516986 410614
rect 517542 410058 552986 410614
rect 553542 410058 591102 410614
rect 591658 410058 592650 410614
rect -8726 410026 592650 410058
rect -6806 406894 590730 406926
rect -6806 406338 -5814 406894
rect -5258 406338 9266 406894
rect 9822 406338 45266 406894
rect 45822 406338 81266 406894
rect 81822 406338 117266 406894
rect 117822 406338 153266 406894
rect 153822 406338 189266 406894
rect 189822 406338 225266 406894
rect 225822 406338 405266 406894
rect 405822 406338 441266 406894
rect 441822 406338 477266 406894
rect 477822 406338 513266 406894
rect 513822 406338 549266 406894
rect 549822 406338 589182 406894
rect 589738 406338 590730 406894
rect -6806 406306 590730 406338
rect -4886 403174 588810 403206
rect -4886 402618 -3894 403174
rect -3338 402618 5546 403174
rect 6102 402618 41546 403174
rect 42102 402618 77546 403174
rect 78102 402618 113546 403174
rect 114102 402618 149546 403174
rect 150102 402618 185546 403174
rect 186102 402618 221546 403174
rect 222102 402618 401546 403174
rect 402102 402618 437546 403174
rect 438102 402618 473546 403174
rect 474102 402618 509546 403174
rect 510102 402618 545546 403174
rect 546102 402618 581546 403174
rect 582102 402618 587262 403174
rect 587818 402618 588810 403174
rect -4886 402586 588810 402618
rect -2966 399454 586890 399486
rect -2966 398898 -1974 399454
rect -1418 398898 1826 399454
rect 2382 398898 37826 399454
rect 38382 398898 73826 399454
rect 74382 398898 109826 399454
rect 110382 398898 145826 399454
rect 146382 398898 181826 399454
rect 182382 398898 217826 399454
rect 218382 399218 239250 399454
rect 239486 399218 269970 399454
rect 270206 399218 300690 399454
rect 300926 399218 331410 399454
rect 331646 399218 362130 399454
rect 362366 399218 397826 399454
rect 218382 399134 397826 399218
rect 218382 398898 239250 399134
rect 239486 398898 269970 399134
rect 270206 398898 300690 399134
rect 300926 398898 331410 399134
rect 331646 398898 362130 399134
rect 362366 398898 397826 399134
rect 398382 398898 433826 399454
rect 434382 398898 469826 399454
rect 470382 398898 505826 399454
rect 506382 398898 541826 399454
rect 542382 398898 577826 399454
rect 578382 398898 585342 399454
rect 585898 398898 586890 399454
rect -2966 398866 586890 398898
rect -8726 392614 592650 392646
rect -8726 392058 -8694 392614
rect -8138 392058 30986 392614
rect 31542 392058 66986 392614
rect 67542 392058 102986 392614
rect 103542 392058 138986 392614
rect 139542 392058 174986 392614
rect 175542 392058 210986 392614
rect 211542 392058 390986 392614
rect 391542 392058 426986 392614
rect 427542 392058 462986 392614
rect 463542 392058 498986 392614
rect 499542 392058 534986 392614
rect 535542 392058 570986 392614
rect 571542 392058 592062 392614
rect 592618 392058 592650 392614
rect -8726 392026 592650 392058
rect -6806 388894 590730 388926
rect -6806 388338 -6774 388894
rect -6218 388338 27266 388894
rect 27822 388338 63266 388894
rect 63822 388338 99266 388894
rect 99822 388338 135266 388894
rect 135822 388338 171266 388894
rect 171822 388338 207266 388894
rect 207822 388338 387266 388894
rect 387822 388338 423266 388894
rect 423822 388338 459266 388894
rect 459822 388338 495266 388894
rect 495822 388338 531266 388894
rect 531822 388338 567266 388894
rect 567822 388338 590142 388894
rect 590698 388338 590730 388894
rect -6806 388306 590730 388338
rect -4886 385174 588810 385206
rect -4886 384618 -4854 385174
rect -4298 384618 23546 385174
rect 24102 384618 59546 385174
rect 60102 384618 95546 385174
rect 96102 384618 131546 385174
rect 132102 384618 167546 385174
rect 168102 384618 203546 385174
rect 204102 384618 419546 385174
rect 420102 384618 455546 385174
rect 456102 384618 491546 385174
rect 492102 384618 527546 385174
rect 528102 384618 563546 385174
rect 564102 384618 588222 385174
rect 588778 384618 588810 385174
rect -4886 384586 588810 384618
rect -2966 381454 586890 381486
rect -2966 380898 -2934 381454
rect -2378 380898 19826 381454
rect 20382 380898 55826 381454
rect 56382 380898 91826 381454
rect 92382 380898 127826 381454
rect 128382 380898 163826 381454
rect 164382 380898 199826 381454
rect 200382 381218 254610 381454
rect 254846 381218 285330 381454
rect 285566 381218 316050 381454
rect 316286 381218 346770 381454
rect 347006 381218 377490 381454
rect 377726 381218 415826 381454
rect 200382 381134 415826 381218
rect 200382 380898 254610 381134
rect 254846 380898 285330 381134
rect 285566 380898 316050 381134
rect 316286 380898 346770 381134
rect 347006 380898 377490 381134
rect 377726 380898 415826 381134
rect 416382 380898 451826 381454
rect 452382 380898 487826 381454
rect 488382 380898 523826 381454
rect 524382 380898 559826 381454
rect 560382 380898 586302 381454
rect 586858 380898 586890 381454
rect -2966 380866 586890 380898
rect -8726 374614 592650 374646
rect -8726 374058 -7734 374614
rect -7178 374058 12986 374614
rect 13542 374058 48986 374614
rect 49542 374058 84986 374614
rect 85542 374058 120986 374614
rect 121542 374058 156986 374614
rect 157542 374058 192986 374614
rect 193542 374058 228986 374614
rect 229542 374058 408986 374614
rect 409542 374058 444986 374614
rect 445542 374058 480986 374614
rect 481542 374058 516986 374614
rect 517542 374058 552986 374614
rect 553542 374058 591102 374614
rect 591658 374058 592650 374614
rect -8726 374026 592650 374058
rect -6806 370894 590730 370926
rect -6806 370338 -5814 370894
rect -5258 370338 9266 370894
rect 9822 370338 45266 370894
rect 45822 370338 81266 370894
rect 81822 370338 117266 370894
rect 117822 370338 153266 370894
rect 153822 370338 189266 370894
rect 189822 370338 225266 370894
rect 225822 370338 405266 370894
rect 405822 370338 441266 370894
rect 441822 370338 477266 370894
rect 477822 370338 513266 370894
rect 513822 370338 549266 370894
rect 549822 370338 589182 370894
rect 589738 370338 590730 370894
rect -6806 370306 590730 370338
rect -4886 367174 588810 367206
rect -4886 366618 -3894 367174
rect -3338 366618 5546 367174
rect 6102 366618 41546 367174
rect 42102 366618 77546 367174
rect 78102 366618 113546 367174
rect 114102 366618 149546 367174
rect 150102 366618 185546 367174
rect 186102 366618 221546 367174
rect 222102 366618 401546 367174
rect 402102 366618 437546 367174
rect 438102 366618 473546 367174
rect 474102 366618 509546 367174
rect 510102 366618 545546 367174
rect 546102 366618 581546 367174
rect 582102 366618 587262 367174
rect 587818 366618 588810 367174
rect -4886 366586 588810 366618
rect -2966 363454 586890 363486
rect -2966 362898 -1974 363454
rect -1418 362898 1826 363454
rect 2382 362898 37826 363454
rect 38382 362898 73826 363454
rect 74382 362898 109826 363454
rect 110382 362898 145826 363454
rect 146382 362898 181826 363454
rect 182382 362898 217826 363454
rect 218382 363218 239250 363454
rect 239486 363218 269970 363454
rect 270206 363218 300690 363454
rect 300926 363218 331410 363454
rect 331646 363218 362130 363454
rect 362366 363218 397826 363454
rect 218382 363134 397826 363218
rect 218382 362898 239250 363134
rect 239486 362898 269970 363134
rect 270206 362898 300690 363134
rect 300926 362898 331410 363134
rect 331646 362898 362130 363134
rect 362366 362898 397826 363134
rect 398382 362898 433826 363454
rect 434382 362898 469826 363454
rect 470382 362898 505826 363454
rect 506382 362898 541826 363454
rect 542382 362898 577826 363454
rect 578382 362898 585342 363454
rect 585898 362898 586890 363454
rect -2966 362866 586890 362898
rect -8726 356614 592650 356646
rect -8726 356058 -8694 356614
rect -8138 356058 30986 356614
rect 31542 356058 66986 356614
rect 67542 356058 102986 356614
rect 103542 356058 138986 356614
rect 139542 356058 174986 356614
rect 175542 356058 210986 356614
rect 211542 356058 390986 356614
rect 391542 356058 426986 356614
rect 427542 356058 462986 356614
rect 463542 356058 498986 356614
rect 499542 356058 534986 356614
rect 535542 356058 570986 356614
rect 571542 356058 592062 356614
rect 592618 356058 592650 356614
rect -8726 356026 592650 356058
rect -6806 352894 590730 352926
rect -6806 352338 -6774 352894
rect -6218 352338 27266 352894
rect 27822 352338 63266 352894
rect 63822 352338 99266 352894
rect 99822 352338 135266 352894
rect 135822 352338 171266 352894
rect 171822 352338 207266 352894
rect 207822 352338 387266 352894
rect 387822 352338 423266 352894
rect 423822 352338 459266 352894
rect 459822 352338 495266 352894
rect 495822 352338 531266 352894
rect 531822 352338 567266 352894
rect 567822 352338 590142 352894
rect 590698 352338 590730 352894
rect -6806 352306 590730 352338
rect -4886 349174 588810 349206
rect -4886 348618 -4854 349174
rect -4298 348618 23546 349174
rect 24102 348618 59546 349174
rect 60102 348618 95546 349174
rect 96102 348618 131546 349174
rect 132102 348618 167546 349174
rect 168102 348618 203546 349174
rect 204102 348618 419546 349174
rect 420102 348618 455546 349174
rect 456102 348618 491546 349174
rect 492102 348618 527546 349174
rect 528102 348618 563546 349174
rect 564102 348618 588222 349174
rect 588778 348618 588810 349174
rect -4886 348586 588810 348618
rect -2966 345454 586890 345486
rect -2966 344898 -2934 345454
rect -2378 344898 19826 345454
rect 20382 344898 55826 345454
rect 56382 344898 91826 345454
rect 92382 344898 127826 345454
rect 128382 344898 163826 345454
rect 164382 344898 199826 345454
rect 200382 345218 254610 345454
rect 254846 345218 285330 345454
rect 285566 345218 316050 345454
rect 316286 345218 346770 345454
rect 347006 345218 377490 345454
rect 377726 345218 415826 345454
rect 200382 345134 415826 345218
rect 200382 344898 254610 345134
rect 254846 344898 285330 345134
rect 285566 344898 316050 345134
rect 316286 344898 346770 345134
rect 347006 344898 377490 345134
rect 377726 344898 415826 345134
rect 416382 344898 451826 345454
rect 452382 344898 487826 345454
rect 488382 344898 523826 345454
rect 524382 344898 559826 345454
rect 560382 344898 586302 345454
rect 586858 344898 586890 345454
rect -2966 344866 586890 344898
rect -8726 338614 592650 338646
rect -8726 338058 -7734 338614
rect -7178 338058 12986 338614
rect 13542 338058 48986 338614
rect 49542 338058 84986 338614
rect 85542 338058 120986 338614
rect 121542 338058 156986 338614
rect 157542 338058 192986 338614
rect 193542 338058 228986 338614
rect 229542 338058 408986 338614
rect 409542 338058 444986 338614
rect 445542 338058 480986 338614
rect 481542 338058 516986 338614
rect 517542 338058 552986 338614
rect 553542 338058 591102 338614
rect 591658 338058 592650 338614
rect -8726 338026 592650 338058
rect -6806 334894 590730 334926
rect -6806 334338 -5814 334894
rect -5258 334338 9266 334894
rect 9822 334338 45266 334894
rect 45822 334338 81266 334894
rect 81822 334338 117266 334894
rect 117822 334338 153266 334894
rect 153822 334338 189266 334894
rect 189822 334338 225266 334894
rect 225822 334338 261266 334894
rect 261822 334338 297266 334894
rect 297822 334338 333266 334894
rect 333822 334338 369266 334894
rect 369822 334338 405266 334894
rect 405822 334338 441266 334894
rect 441822 334338 477266 334894
rect 477822 334338 513266 334894
rect 513822 334338 549266 334894
rect 549822 334338 589182 334894
rect 589738 334338 590730 334894
rect -6806 334306 590730 334338
rect -4886 331174 588810 331206
rect -4886 330618 -3894 331174
rect -3338 330618 5546 331174
rect 6102 330618 41546 331174
rect 42102 330618 77546 331174
rect 78102 330618 113546 331174
rect 114102 330618 149546 331174
rect 150102 330618 185546 331174
rect 186102 330618 221546 331174
rect 222102 330618 257546 331174
rect 258102 330618 293546 331174
rect 294102 330618 329546 331174
rect 330102 330618 365546 331174
rect 366102 330618 401546 331174
rect 402102 330618 437546 331174
rect 438102 330618 473546 331174
rect 474102 330618 509546 331174
rect 510102 330618 545546 331174
rect 546102 330618 581546 331174
rect 582102 330618 587262 331174
rect 587818 330618 588810 331174
rect -4886 330586 588810 330618
rect -2966 327454 586890 327486
rect -2966 326898 -1974 327454
rect -1418 326898 1826 327454
rect 2382 326898 37826 327454
rect 38382 326898 73826 327454
rect 74382 326898 109826 327454
rect 110382 326898 145826 327454
rect 146382 326898 181826 327454
rect 182382 326898 217826 327454
rect 218382 326898 253826 327454
rect 254382 326898 289826 327454
rect 290382 326898 325826 327454
rect 326382 326898 361826 327454
rect 362382 326898 397826 327454
rect 398382 326898 433826 327454
rect 434382 326898 469826 327454
rect 470382 326898 505826 327454
rect 506382 326898 541826 327454
rect 542382 326898 577826 327454
rect 578382 326898 585342 327454
rect 585898 326898 586890 327454
rect -2966 326866 586890 326898
rect -8726 320614 592650 320646
rect -8726 320058 -8694 320614
rect -8138 320058 30986 320614
rect 31542 320058 66986 320614
rect 67542 320058 102986 320614
rect 103542 320058 138986 320614
rect 139542 320058 174986 320614
rect 175542 320058 210986 320614
rect 211542 320058 246986 320614
rect 247542 320058 282986 320614
rect 283542 320058 318986 320614
rect 319542 320058 354986 320614
rect 355542 320058 390986 320614
rect 391542 320058 426986 320614
rect 427542 320058 462986 320614
rect 463542 320058 498986 320614
rect 499542 320058 534986 320614
rect 535542 320058 570986 320614
rect 571542 320058 592062 320614
rect 592618 320058 592650 320614
rect -8726 320026 592650 320058
rect -6806 316894 590730 316926
rect -6806 316338 -6774 316894
rect -6218 316338 27266 316894
rect 27822 316338 63266 316894
rect 63822 316338 99266 316894
rect 99822 316338 135266 316894
rect 135822 316338 171266 316894
rect 171822 316338 207266 316894
rect 207822 316338 243266 316894
rect 243822 316338 279266 316894
rect 279822 316338 315266 316894
rect 315822 316338 351266 316894
rect 351822 316338 387266 316894
rect 387822 316338 423266 316894
rect 423822 316338 459266 316894
rect 459822 316338 495266 316894
rect 495822 316338 531266 316894
rect 531822 316338 567266 316894
rect 567822 316338 590142 316894
rect 590698 316338 590730 316894
rect -6806 316306 590730 316338
rect -4886 313174 588810 313206
rect -4886 312618 -4854 313174
rect -4298 312618 23546 313174
rect 24102 312618 59546 313174
rect 60102 312618 95546 313174
rect 96102 312618 131546 313174
rect 132102 312618 167546 313174
rect 168102 312618 203546 313174
rect 204102 312618 239546 313174
rect 240102 312618 275546 313174
rect 276102 312618 311546 313174
rect 312102 312618 347546 313174
rect 348102 312618 383546 313174
rect 384102 312618 419546 313174
rect 420102 312618 455546 313174
rect 456102 312618 491546 313174
rect 492102 312618 527546 313174
rect 528102 312618 563546 313174
rect 564102 312618 588222 313174
rect 588778 312618 588810 313174
rect -4886 312586 588810 312618
rect -2966 309454 586890 309486
rect -2966 308898 -2934 309454
rect -2378 308898 19826 309454
rect 20382 308898 55826 309454
rect 56382 308898 91826 309454
rect 92382 308898 127826 309454
rect 128382 308898 163826 309454
rect 164382 308898 199826 309454
rect 200382 308898 235826 309454
rect 236382 308898 271826 309454
rect 272382 308898 307826 309454
rect 308382 308898 343826 309454
rect 344382 308898 379826 309454
rect 380382 308898 415826 309454
rect 416382 308898 451826 309454
rect 452382 308898 487826 309454
rect 488382 308898 523826 309454
rect 524382 308898 559826 309454
rect 560382 308898 586302 309454
rect 586858 308898 586890 309454
rect -2966 308866 586890 308898
rect -8726 302614 592650 302646
rect -8726 302058 -7734 302614
rect -7178 302058 12986 302614
rect 13542 302058 48986 302614
rect 49542 302058 84986 302614
rect 85542 302058 120986 302614
rect 121542 302058 156986 302614
rect 157542 302058 192986 302614
rect 193542 302058 228986 302614
rect 229542 302058 264986 302614
rect 265542 302058 300986 302614
rect 301542 302058 336986 302614
rect 337542 302058 372986 302614
rect 373542 302058 408986 302614
rect 409542 302058 444986 302614
rect 445542 302058 480986 302614
rect 481542 302058 516986 302614
rect 517542 302058 552986 302614
rect 553542 302058 591102 302614
rect 591658 302058 592650 302614
rect -8726 302026 592650 302058
rect -6806 298894 590730 298926
rect -6806 298338 -5814 298894
rect -5258 298338 9266 298894
rect 9822 298338 45266 298894
rect 45822 298338 81266 298894
rect 81822 298338 117266 298894
rect 117822 298338 153266 298894
rect 153822 298338 189266 298894
rect 189822 298338 225266 298894
rect 225822 298338 261266 298894
rect 261822 298338 297266 298894
rect 297822 298338 333266 298894
rect 333822 298338 369266 298894
rect 369822 298338 405266 298894
rect 405822 298338 441266 298894
rect 441822 298338 477266 298894
rect 477822 298338 513266 298894
rect 513822 298338 549266 298894
rect 549822 298338 589182 298894
rect 589738 298338 590730 298894
rect -6806 298306 590730 298338
rect -4886 295174 588810 295206
rect -4886 294618 -3894 295174
rect -3338 294618 5546 295174
rect 6102 294618 41546 295174
rect 42102 294618 77546 295174
rect 78102 294618 113546 295174
rect 114102 294618 149546 295174
rect 150102 294618 185546 295174
rect 186102 294618 221546 295174
rect 222102 294618 257546 295174
rect 258102 294618 293546 295174
rect 294102 294618 329546 295174
rect 330102 294618 365546 295174
rect 366102 294618 401546 295174
rect 402102 294618 437546 295174
rect 438102 294618 473546 295174
rect 474102 294618 509546 295174
rect 510102 294618 545546 295174
rect 546102 294618 581546 295174
rect 582102 294618 587262 295174
rect 587818 294618 588810 295174
rect -4886 294586 588810 294618
rect -2966 291454 586890 291486
rect -2966 290898 -1974 291454
rect -1418 290898 1826 291454
rect 2382 290898 37826 291454
rect 38382 290898 73826 291454
rect 74382 290898 109826 291454
rect 110382 290898 145826 291454
rect 146382 290898 181826 291454
rect 182382 290898 217826 291454
rect 218382 290898 253826 291454
rect 254382 290898 289826 291454
rect 290382 290898 325826 291454
rect 326382 290898 361826 291454
rect 362382 290898 397826 291454
rect 398382 290898 433826 291454
rect 434382 290898 469826 291454
rect 470382 290898 505826 291454
rect 506382 290898 541826 291454
rect 542382 290898 577826 291454
rect 578382 290898 585342 291454
rect 585898 290898 586890 291454
rect -2966 290866 586890 290898
rect -8726 284614 592650 284646
rect -8726 284058 -8694 284614
rect -8138 284058 30986 284614
rect 31542 284058 66986 284614
rect 67542 284058 102986 284614
rect 103542 284058 138986 284614
rect 139542 284058 174986 284614
rect 175542 284058 210986 284614
rect 211542 284058 246986 284614
rect 247542 284058 282986 284614
rect 283542 284058 318986 284614
rect 319542 284058 354986 284614
rect 355542 284058 390986 284614
rect 391542 284058 426986 284614
rect 427542 284058 462986 284614
rect 463542 284058 498986 284614
rect 499542 284058 534986 284614
rect 535542 284058 570986 284614
rect 571542 284058 592062 284614
rect 592618 284058 592650 284614
rect -8726 284026 592650 284058
rect -6806 280894 590730 280926
rect -6806 280338 -6774 280894
rect -6218 280338 27266 280894
rect 27822 280338 63266 280894
rect 63822 280338 99266 280894
rect 99822 280338 135266 280894
rect 135822 280338 171266 280894
rect 171822 280338 207266 280894
rect 207822 280338 243266 280894
rect 243822 280338 279266 280894
rect 279822 280338 315266 280894
rect 315822 280338 351266 280894
rect 351822 280338 387266 280894
rect 387822 280338 423266 280894
rect 423822 280338 459266 280894
rect 459822 280338 495266 280894
rect 495822 280338 531266 280894
rect 531822 280338 567266 280894
rect 567822 280338 590142 280894
rect 590698 280338 590730 280894
rect -6806 280306 590730 280338
rect -4886 277174 588810 277206
rect -4886 276618 -4854 277174
rect -4298 276618 23546 277174
rect 24102 276618 59546 277174
rect 60102 276618 95546 277174
rect 96102 276618 131546 277174
rect 132102 276618 167546 277174
rect 168102 276618 203546 277174
rect 204102 276618 239546 277174
rect 240102 276618 275546 277174
rect 276102 276618 311546 277174
rect 312102 276618 347546 277174
rect 348102 276618 383546 277174
rect 384102 276618 419546 277174
rect 420102 276618 455546 277174
rect 456102 276618 491546 277174
rect 492102 276618 527546 277174
rect 528102 276618 563546 277174
rect 564102 276618 588222 277174
rect 588778 276618 588810 277174
rect -4886 276586 588810 276618
rect -2966 273454 586890 273486
rect -2966 272898 -2934 273454
rect -2378 272898 19826 273454
rect 20382 272898 55826 273454
rect 56382 272898 91826 273454
rect 92382 272898 127826 273454
rect 128382 272898 163826 273454
rect 164382 272898 199826 273454
rect 200382 272898 235826 273454
rect 236382 272898 271826 273454
rect 272382 272898 307826 273454
rect 308382 272898 343826 273454
rect 344382 272898 379826 273454
rect 380382 272898 415826 273454
rect 416382 272898 451826 273454
rect 452382 272898 487826 273454
rect 488382 272898 523826 273454
rect 524382 272898 559826 273454
rect 560382 272898 586302 273454
rect 586858 272898 586890 273454
rect -2966 272866 586890 272898
rect -8726 266614 592650 266646
rect -8726 266058 -7734 266614
rect -7178 266058 12986 266614
rect 13542 266058 48986 266614
rect 49542 266058 84986 266614
rect 85542 266058 120986 266614
rect 121542 266058 156986 266614
rect 157542 266058 192986 266614
rect 193542 266058 228986 266614
rect 229542 266058 264986 266614
rect 265542 266058 300986 266614
rect 301542 266058 336986 266614
rect 337542 266058 372986 266614
rect 373542 266058 408986 266614
rect 409542 266058 444986 266614
rect 445542 266058 480986 266614
rect 481542 266058 516986 266614
rect 517542 266058 552986 266614
rect 553542 266058 591102 266614
rect 591658 266058 592650 266614
rect -8726 266026 592650 266058
rect -6806 262894 590730 262926
rect -6806 262338 -5814 262894
rect -5258 262338 9266 262894
rect 9822 262338 45266 262894
rect 45822 262338 81266 262894
rect 81822 262338 117266 262894
rect 117822 262338 153266 262894
rect 153822 262338 189266 262894
rect 189822 262338 225266 262894
rect 225822 262338 261266 262894
rect 261822 262338 297266 262894
rect 297822 262338 333266 262894
rect 333822 262338 369266 262894
rect 369822 262338 405266 262894
rect 405822 262338 441266 262894
rect 441822 262338 477266 262894
rect 477822 262338 513266 262894
rect 513822 262338 549266 262894
rect 549822 262338 589182 262894
rect 589738 262338 590730 262894
rect -6806 262306 590730 262338
rect -4886 259174 588810 259206
rect -4886 258618 -3894 259174
rect -3338 258618 5546 259174
rect 6102 258618 41546 259174
rect 42102 258618 77546 259174
rect 78102 258618 113546 259174
rect 114102 258618 149546 259174
rect 150102 258618 185546 259174
rect 186102 258618 221546 259174
rect 222102 258618 257546 259174
rect 258102 258618 293546 259174
rect 294102 258618 329546 259174
rect 330102 258618 365546 259174
rect 366102 258618 401546 259174
rect 402102 258618 437546 259174
rect 438102 258618 473546 259174
rect 474102 258618 509546 259174
rect 510102 258618 545546 259174
rect 546102 258618 581546 259174
rect 582102 258618 587262 259174
rect 587818 258618 588810 259174
rect -4886 258586 588810 258618
rect -2966 255454 586890 255486
rect -2966 254898 -1974 255454
rect -1418 254898 1826 255454
rect 2382 254898 37826 255454
rect 38382 254898 73826 255454
rect 74382 254898 109826 255454
rect 110382 254898 145826 255454
rect 146382 254898 181826 255454
rect 182382 254898 217826 255454
rect 218382 254898 253826 255454
rect 254382 254898 289826 255454
rect 290382 254898 325826 255454
rect 326382 254898 361826 255454
rect 362382 254898 397826 255454
rect 398382 254898 433826 255454
rect 434382 254898 469826 255454
rect 470382 254898 505826 255454
rect 506382 254898 541826 255454
rect 542382 254898 577826 255454
rect 578382 254898 585342 255454
rect 585898 254898 586890 255454
rect -2966 254866 586890 254898
rect -8726 248614 592650 248646
rect -8726 248058 -8694 248614
rect -8138 248058 30986 248614
rect 31542 248058 66986 248614
rect 67542 248058 102986 248614
rect 103542 248058 138986 248614
rect 139542 248058 174986 248614
rect 175542 248058 210986 248614
rect 211542 248058 246986 248614
rect 247542 248058 282986 248614
rect 283542 248058 318986 248614
rect 319542 248058 354986 248614
rect 355542 248058 390986 248614
rect 391542 248058 426986 248614
rect 427542 248058 462986 248614
rect 463542 248058 498986 248614
rect 499542 248058 534986 248614
rect 535542 248058 570986 248614
rect 571542 248058 592062 248614
rect 592618 248058 592650 248614
rect -8726 248026 592650 248058
rect -6806 244894 590730 244926
rect -6806 244338 -6774 244894
rect -6218 244338 27266 244894
rect 27822 244338 63266 244894
rect 63822 244338 99266 244894
rect 99822 244338 135266 244894
rect 135822 244338 171266 244894
rect 171822 244338 207266 244894
rect 207822 244338 243266 244894
rect 243822 244338 279266 244894
rect 279822 244338 315266 244894
rect 315822 244338 351266 244894
rect 351822 244338 387266 244894
rect 387822 244338 423266 244894
rect 423822 244338 459266 244894
rect 459822 244338 495266 244894
rect 495822 244338 531266 244894
rect 531822 244338 567266 244894
rect 567822 244338 590142 244894
rect 590698 244338 590730 244894
rect -6806 244306 590730 244338
rect -4886 241174 588810 241206
rect -4886 240618 -4854 241174
rect -4298 240618 23546 241174
rect 24102 240618 59546 241174
rect 60102 240618 95546 241174
rect 96102 240618 131546 241174
rect 132102 240618 167546 241174
rect 168102 240618 203546 241174
rect 204102 240618 239546 241174
rect 240102 240618 275546 241174
rect 276102 240618 311546 241174
rect 312102 240618 347546 241174
rect 348102 240618 383546 241174
rect 384102 240618 419546 241174
rect 420102 240618 455546 241174
rect 456102 240618 491546 241174
rect 492102 240618 527546 241174
rect 528102 240618 563546 241174
rect 564102 240618 588222 241174
rect 588778 240618 588810 241174
rect -4886 240586 588810 240618
rect -2966 237454 586890 237486
rect -2966 236898 -2934 237454
rect -2378 236898 19826 237454
rect 20382 236898 55826 237454
rect 56382 236898 91826 237454
rect 92382 236898 127826 237454
rect 128382 236898 163826 237454
rect 164382 236898 199826 237454
rect 200382 236898 235826 237454
rect 236382 236898 271826 237454
rect 272382 236898 307826 237454
rect 308382 236898 343826 237454
rect 344382 236898 379826 237454
rect 380382 236898 415826 237454
rect 416382 236898 451826 237454
rect 452382 236898 487826 237454
rect 488382 236898 523826 237454
rect 524382 236898 559826 237454
rect 560382 236898 586302 237454
rect 586858 236898 586890 237454
rect -2966 236866 586890 236898
rect -8726 230614 592650 230646
rect -8726 230058 -7734 230614
rect -7178 230058 12986 230614
rect 13542 230058 48986 230614
rect 49542 230058 84986 230614
rect 85542 230058 120986 230614
rect 121542 230058 156986 230614
rect 157542 230058 192986 230614
rect 193542 230058 228986 230614
rect 229542 230058 264986 230614
rect 265542 230058 300986 230614
rect 301542 230058 336986 230614
rect 337542 230058 372986 230614
rect 373542 230058 408986 230614
rect 409542 230058 444986 230614
rect 445542 230058 480986 230614
rect 481542 230058 516986 230614
rect 517542 230058 552986 230614
rect 553542 230058 591102 230614
rect 591658 230058 592650 230614
rect -8726 230026 592650 230058
rect -6806 226894 590730 226926
rect -6806 226338 -5814 226894
rect -5258 226338 9266 226894
rect 9822 226338 45266 226894
rect 45822 226338 81266 226894
rect 81822 226338 117266 226894
rect 117822 226338 153266 226894
rect 153822 226338 189266 226894
rect 189822 226338 225266 226894
rect 225822 226338 261266 226894
rect 261822 226338 297266 226894
rect 297822 226338 333266 226894
rect 333822 226338 369266 226894
rect 369822 226338 405266 226894
rect 405822 226338 441266 226894
rect 441822 226338 477266 226894
rect 477822 226338 513266 226894
rect 513822 226338 549266 226894
rect 549822 226338 589182 226894
rect 589738 226338 590730 226894
rect -6806 226306 590730 226338
rect -4886 223174 588810 223206
rect -4886 222618 -3894 223174
rect -3338 222618 5546 223174
rect 6102 222618 41546 223174
rect 42102 222618 77546 223174
rect 78102 222618 113546 223174
rect 114102 222618 149546 223174
rect 150102 222618 185546 223174
rect 186102 222618 221546 223174
rect 222102 222618 257546 223174
rect 258102 222618 293546 223174
rect 294102 222618 329546 223174
rect 330102 222618 365546 223174
rect 366102 222618 401546 223174
rect 402102 222618 437546 223174
rect 438102 222618 473546 223174
rect 474102 222618 509546 223174
rect 510102 222618 545546 223174
rect 546102 222618 581546 223174
rect 582102 222618 587262 223174
rect 587818 222618 588810 223174
rect -4886 222586 588810 222618
rect -2966 219454 586890 219486
rect -2966 218898 -1974 219454
rect -1418 218898 1826 219454
rect 2382 218898 37826 219454
rect 38382 218898 73826 219454
rect 74382 218898 109826 219454
rect 110382 218898 145826 219454
rect 146382 218898 181826 219454
rect 182382 218898 217826 219454
rect 218382 218898 253826 219454
rect 254382 218898 289826 219454
rect 290382 218898 325826 219454
rect 326382 218898 361826 219454
rect 362382 218898 397826 219454
rect 398382 218898 433826 219454
rect 434382 218898 469826 219454
rect 470382 218898 505826 219454
rect 506382 218898 541826 219454
rect 542382 218898 577826 219454
rect 578382 218898 585342 219454
rect 585898 218898 586890 219454
rect -2966 218866 586890 218898
rect -8726 212614 592650 212646
rect -8726 212058 -8694 212614
rect -8138 212058 30986 212614
rect 31542 212058 66986 212614
rect 67542 212058 102986 212614
rect 103542 212058 138986 212614
rect 139542 212058 174986 212614
rect 175542 212058 210986 212614
rect 211542 212058 246986 212614
rect 247542 212058 282986 212614
rect 283542 212058 318986 212614
rect 319542 212058 354986 212614
rect 355542 212058 390986 212614
rect 391542 212058 426986 212614
rect 427542 212058 462986 212614
rect 463542 212058 498986 212614
rect 499542 212058 534986 212614
rect 535542 212058 570986 212614
rect 571542 212058 592062 212614
rect 592618 212058 592650 212614
rect -8726 212026 592650 212058
rect -6806 208894 590730 208926
rect -6806 208338 -6774 208894
rect -6218 208338 27266 208894
rect 27822 208338 63266 208894
rect 63822 208338 99266 208894
rect 99822 208338 135266 208894
rect 135822 208338 171266 208894
rect 171822 208338 207266 208894
rect 207822 208338 243266 208894
rect 243822 208338 279266 208894
rect 279822 208338 315266 208894
rect 315822 208338 351266 208894
rect 351822 208338 387266 208894
rect 387822 208338 423266 208894
rect 423822 208338 459266 208894
rect 459822 208338 495266 208894
rect 495822 208338 531266 208894
rect 531822 208338 567266 208894
rect 567822 208338 590142 208894
rect 590698 208338 590730 208894
rect -6806 208306 590730 208338
rect -4886 205174 588810 205206
rect -4886 204618 -4854 205174
rect -4298 204618 23546 205174
rect 24102 204618 59546 205174
rect 60102 204618 95546 205174
rect 96102 204618 131546 205174
rect 132102 204618 167546 205174
rect 168102 204618 203546 205174
rect 204102 204618 239546 205174
rect 240102 204618 275546 205174
rect 276102 204618 311546 205174
rect 312102 204618 347546 205174
rect 348102 204618 383546 205174
rect 384102 204618 419546 205174
rect 420102 204618 455546 205174
rect 456102 204618 491546 205174
rect 492102 204618 527546 205174
rect 528102 204618 563546 205174
rect 564102 204618 588222 205174
rect 588778 204618 588810 205174
rect -4886 204586 588810 204618
rect -2966 201454 586890 201486
rect -2966 200898 -2934 201454
rect -2378 200898 19826 201454
rect 20382 200898 55826 201454
rect 56382 200898 91826 201454
rect 92382 200898 127826 201454
rect 128382 200898 163826 201454
rect 164382 200898 199826 201454
rect 200382 200898 235826 201454
rect 236382 200898 271826 201454
rect 272382 200898 307826 201454
rect 308382 200898 343826 201454
rect 344382 200898 379826 201454
rect 380382 200898 415826 201454
rect 416382 200898 451826 201454
rect 452382 200898 487826 201454
rect 488382 200898 523826 201454
rect 524382 200898 559826 201454
rect 560382 200898 586302 201454
rect 586858 200898 586890 201454
rect -2966 200866 586890 200898
rect -8726 194614 592650 194646
rect -8726 194058 -7734 194614
rect -7178 194058 12986 194614
rect 13542 194058 48986 194614
rect 49542 194058 84986 194614
rect 85542 194058 120986 194614
rect 121542 194058 156986 194614
rect 157542 194058 192986 194614
rect 193542 194058 228986 194614
rect 229542 194058 264986 194614
rect 265542 194058 300986 194614
rect 301542 194058 336986 194614
rect 337542 194058 372986 194614
rect 373542 194058 408986 194614
rect 409542 194058 444986 194614
rect 445542 194058 480986 194614
rect 481542 194058 516986 194614
rect 517542 194058 552986 194614
rect 553542 194058 591102 194614
rect 591658 194058 592650 194614
rect -8726 194026 592650 194058
rect -6806 190894 590730 190926
rect -6806 190338 -5814 190894
rect -5258 190338 9266 190894
rect 9822 190338 45266 190894
rect 45822 190338 81266 190894
rect 81822 190338 117266 190894
rect 117822 190338 153266 190894
rect 153822 190338 189266 190894
rect 189822 190338 225266 190894
rect 225822 190338 261266 190894
rect 261822 190338 297266 190894
rect 297822 190338 333266 190894
rect 333822 190338 369266 190894
rect 369822 190338 405266 190894
rect 405822 190338 441266 190894
rect 441822 190338 477266 190894
rect 477822 190338 513266 190894
rect 513822 190338 549266 190894
rect 549822 190338 589182 190894
rect 589738 190338 590730 190894
rect -6806 190306 590730 190338
rect -4886 187174 588810 187206
rect -4886 186618 -3894 187174
rect -3338 186618 5546 187174
rect 6102 186618 41546 187174
rect 42102 186618 77546 187174
rect 78102 186618 113546 187174
rect 114102 186618 149546 187174
rect 150102 186618 185546 187174
rect 186102 186618 221546 187174
rect 222102 186618 257546 187174
rect 258102 186618 293546 187174
rect 294102 186618 329546 187174
rect 330102 186618 365546 187174
rect 366102 186618 401546 187174
rect 402102 186618 437546 187174
rect 438102 186618 473546 187174
rect 474102 186618 509546 187174
rect 510102 186618 545546 187174
rect 546102 186618 581546 187174
rect 582102 186618 587262 187174
rect 587818 186618 588810 187174
rect -4886 186586 588810 186618
rect -2966 183454 586890 183486
rect -2966 182898 -1974 183454
rect -1418 182898 1826 183454
rect 2382 182898 37826 183454
rect 38382 182898 73826 183454
rect 74382 182898 109826 183454
rect 110382 182898 145826 183454
rect 146382 182898 181826 183454
rect 182382 182898 217826 183454
rect 218382 182898 253826 183454
rect 254382 182898 289826 183454
rect 290382 182898 325826 183454
rect 326382 182898 361826 183454
rect 362382 182898 397826 183454
rect 398382 182898 433826 183454
rect 434382 182898 469826 183454
rect 470382 182898 505826 183454
rect 506382 182898 541826 183454
rect 542382 182898 577826 183454
rect 578382 182898 585342 183454
rect 585898 182898 586890 183454
rect -2966 182866 586890 182898
rect -8726 176614 592650 176646
rect -8726 176058 -8694 176614
rect -8138 176058 30986 176614
rect 31542 176058 66986 176614
rect 67542 176058 102986 176614
rect 103542 176058 138986 176614
rect 139542 176058 174986 176614
rect 175542 176058 210986 176614
rect 211542 176058 246986 176614
rect 247542 176058 282986 176614
rect 283542 176058 318986 176614
rect 319542 176058 354986 176614
rect 355542 176058 390986 176614
rect 391542 176058 426986 176614
rect 427542 176058 462986 176614
rect 463542 176058 498986 176614
rect 499542 176058 534986 176614
rect 535542 176058 570986 176614
rect 571542 176058 592062 176614
rect 592618 176058 592650 176614
rect -8726 176026 592650 176058
rect -6806 172894 590730 172926
rect -6806 172338 -6774 172894
rect -6218 172338 27266 172894
rect 27822 172338 63266 172894
rect 63822 172338 99266 172894
rect 99822 172338 135266 172894
rect 135822 172338 171266 172894
rect 171822 172338 207266 172894
rect 207822 172338 243266 172894
rect 243822 172338 279266 172894
rect 279822 172338 315266 172894
rect 315822 172338 351266 172894
rect 351822 172338 387266 172894
rect 387822 172338 423266 172894
rect 423822 172338 459266 172894
rect 459822 172338 495266 172894
rect 495822 172338 531266 172894
rect 531822 172338 567266 172894
rect 567822 172338 590142 172894
rect 590698 172338 590730 172894
rect -6806 172306 590730 172338
rect -4886 169174 588810 169206
rect -4886 168618 -4854 169174
rect -4298 168618 23546 169174
rect 24102 168618 59546 169174
rect 60102 168618 95546 169174
rect 96102 168618 131546 169174
rect 132102 168618 167546 169174
rect 168102 168618 203546 169174
rect 204102 168618 239546 169174
rect 240102 168618 275546 169174
rect 276102 168618 311546 169174
rect 312102 168618 347546 169174
rect 348102 168618 383546 169174
rect 384102 168618 419546 169174
rect 420102 168618 455546 169174
rect 456102 168618 491546 169174
rect 492102 168618 527546 169174
rect 528102 168618 563546 169174
rect 564102 168618 588222 169174
rect 588778 168618 588810 169174
rect -4886 168586 588810 168618
rect -2966 165454 586890 165486
rect -2966 164898 -2934 165454
rect -2378 164898 19826 165454
rect 20382 164898 55826 165454
rect 56382 164898 91826 165454
rect 92382 164898 127826 165454
rect 128382 164898 163826 165454
rect 164382 164898 199826 165454
rect 200382 164898 235826 165454
rect 236382 164898 271826 165454
rect 272382 164898 307826 165454
rect 308382 164898 343826 165454
rect 344382 164898 379826 165454
rect 380382 164898 415826 165454
rect 416382 164898 451826 165454
rect 452382 164898 487826 165454
rect 488382 164898 523826 165454
rect 524382 164898 559826 165454
rect 560382 164898 586302 165454
rect 586858 164898 586890 165454
rect -2966 164866 586890 164898
rect -8726 158614 592650 158646
rect -8726 158058 -7734 158614
rect -7178 158058 12986 158614
rect 13542 158058 48986 158614
rect 49542 158058 84986 158614
rect 85542 158058 120986 158614
rect 121542 158058 156986 158614
rect 157542 158058 192986 158614
rect 193542 158058 228986 158614
rect 229542 158058 264986 158614
rect 265542 158058 300986 158614
rect 301542 158058 336986 158614
rect 337542 158058 372986 158614
rect 373542 158058 408986 158614
rect 409542 158058 444986 158614
rect 445542 158058 480986 158614
rect 481542 158058 516986 158614
rect 517542 158058 552986 158614
rect 553542 158058 591102 158614
rect 591658 158058 592650 158614
rect -8726 158026 592650 158058
rect -6806 154894 590730 154926
rect -6806 154338 -5814 154894
rect -5258 154338 9266 154894
rect 9822 154338 45266 154894
rect 45822 154338 81266 154894
rect 81822 154338 117266 154894
rect 117822 154338 153266 154894
rect 153822 154338 189266 154894
rect 189822 154338 225266 154894
rect 225822 154338 261266 154894
rect 261822 154338 297266 154894
rect 297822 154338 333266 154894
rect 333822 154338 369266 154894
rect 369822 154338 405266 154894
rect 405822 154338 441266 154894
rect 441822 154338 477266 154894
rect 477822 154338 513266 154894
rect 513822 154338 549266 154894
rect 549822 154338 589182 154894
rect 589738 154338 590730 154894
rect -6806 154306 590730 154338
rect -4886 151174 588810 151206
rect -4886 150618 -3894 151174
rect -3338 150618 5546 151174
rect 6102 150618 41546 151174
rect 42102 150618 77546 151174
rect 78102 150618 113546 151174
rect 114102 150618 149546 151174
rect 150102 150618 185546 151174
rect 186102 150618 221546 151174
rect 222102 150618 257546 151174
rect 258102 150618 293546 151174
rect 294102 150618 329546 151174
rect 330102 150618 365546 151174
rect 366102 150618 401546 151174
rect 402102 150618 437546 151174
rect 438102 150618 473546 151174
rect 474102 150618 509546 151174
rect 510102 150618 545546 151174
rect 546102 150618 581546 151174
rect 582102 150618 587262 151174
rect 587818 150618 588810 151174
rect -4886 150586 588810 150618
rect -2966 147454 586890 147486
rect -2966 146898 -1974 147454
rect -1418 146898 1826 147454
rect 2382 146898 37826 147454
rect 38382 146898 73826 147454
rect 74382 146898 109826 147454
rect 110382 146898 145826 147454
rect 146382 146898 181826 147454
rect 182382 146898 217826 147454
rect 218382 146898 253826 147454
rect 254382 146898 289826 147454
rect 290382 146898 325826 147454
rect 326382 146898 361826 147454
rect 362382 146898 397826 147454
rect 398382 146898 433826 147454
rect 434382 146898 469826 147454
rect 470382 146898 505826 147454
rect 506382 146898 541826 147454
rect 542382 146898 577826 147454
rect 578382 146898 585342 147454
rect 585898 146898 586890 147454
rect -2966 146866 586890 146898
rect -8726 140614 592650 140646
rect -8726 140058 -8694 140614
rect -8138 140058 30986 140614
rect 31542 140058 66986 140614
rect 67542 140058 102986 140614
rect 103542 140058 138986 140614
rect 139542 140058 174986 140614
rect 175542 140058 210986 140614
rect 211542 140058 246986 140614
rect 247542 140058 282986 140614
rect 283542 140058 318986 140614
rect 319542 140058 354986 140614
rect 355542 140058 390986 140614
rect 391542 140058 426986 140614
rect 427542 140058 462986 140614
rect 463542 140058 498986 140614
rect 499542 140058 534986 140614
rect 535542 140058 570986 140614
rect 571542 140058 592062 140614
rect 592618 140058 592650 140614
rect -8726 140026 592650 140058
rect -6806 136894 590730 136926
rect -6806 136338 -6774 136894
rect -6218 136338 27266 136894
rect 27822 136338 63266 136894
rect 63822 136338 99266 136894
rect 99822 136338 135266 136894
rect 135822 136338 171266 136894
rect 171822 136338 207266 136894
rect 207822 136338 243266 136894
rect 243822 136338 279266 136894
rect 279822 136338 315266 136894
rect 315822 136338 351266 136894
rect 351822 136338 387266 136894
rect 387822 136338 423266 136894
rect 423822 136338 459266 136894
rect 459822 136338 495266 136894
rect 495822 136338 531266 136894
rect 531822 136338 567266 136894
rect 567822 136338 590142 136894
rect 590698 136338 590730 136894
rect -6806 136306 590730 136338
rect -4886 133174 588810 133206
rect -4886 132618 -4854 133174
rect -4298 132618 23546 133174
rect 24102 132618 59546 133174
rect 60102 132618 95546 133174
rect 96102 132618 131546 133174
rect 132102 132618 167546 133174
rect 168102 132618 203546 133174
rect 204102 132618 239546 133174
rect 240102 132618 275546 133174
rect 276102 132618 311546 133174
rect 312102 132618 347546 133174
rect 348102 132618 383546 133174
rect 384102 132618 419546 133174
rect 420102 132618 455546 133174
rect 456102 132618 491546 133174
rect 492102 132618 527546 133174
rect 528102 132618 563546 133174
rect 564102 132618 588222 133174
rect 588778 132618 588810 133174
rect -4886 132586 588810 132618
rect -2966 129454 586890 129486
rect -2966 128898 -2934 129454
rect -2378 128898 19826 129454
rect 20382 128898 55826 129454
rect 56382 128898 91826 129454
rect 92382 128898 127826 129454
rect 128382 128898 163826 129454
rect 164382 128898 199826 129454
rect 200382 128898 235826 129454
rect 236382 128898 271826 129454
rect 272382 128898 307826 129454
rect 308382 128898 343826 129454
rect 344382 128898 379826 129454
rect 380382 128898 415826 129454
rect 416382 128898 451826 129454
rect 452382 128898 487826 129454
rect 488382 128898 523826 129454
rect 524382 128898 559826 129454
rect 560382 128898 586302 129454
rect 586858 128898 586890 129454
rect -2966 128866 586890 128898
rect -8726 122614 592650 122646
rect -8726 122058 -7734 122614
rect -7178 122058 12986 122614
rect 13542 122058 48986 122614
rect 49542 122058 84986 122614
rect 85542 122058 120986 122614
rect 121542 122058 156986 122614
rect 157542 122058 192986 122614
rect 193542 122058 228986 122614
rect 229542 122058 264986 122614
rect 265542 122058 300986 122614
rect 301542 122058 336986 122614
rect 337542 122058 372986 122614
rect 373542 122058 408986 122614
rect 409542 122058 444986 122614
rect 445542 122058 480986 122614
rect 481542 122058 516986 122614
rect 517542 122058 552986 122614
rect 553542 122058 591102 122614
rect 591658 122058 592650 122614
rect -8726 122026 592650 122058
rect -6806 118894 590730 118926
rect -6806 118338 -5814 118894
rect -5258 118338 9266 118894
rect 9822 118338 45266 118894
rect 45822 118338 81266 118894
rect 81822 118338 117266 118894
rect 117822 118338 153266 118894
rect 153822 118338 189266 118894
rect 189822 118338 225266 118894
rect 225822 118338 261266 118894
rect 261822 118338 297266 118894
rect 297822 118338 333266 118894
rect 333822 118338 369266 118894
rect 369822 118338 405266 118894
rect 405822 118338 441266 118894
rect 441822 118338 477266 118894
rect 477822 118338 513266 118894
rect 513822 118338 549266 118894
rect 549822 118338 589182 118894
rect 589738 118338 590730 118894
rect -6806 118306 590730 118338
rect -4886 115174 588810 115206
rect -4886 114618 -3894 115174
rect -3338 114618 5546 115174
rect 6102 114618 41546 115174
rect 42102 114618 77546 115174
rect 78102 114618 113546 115174
rect 114102 114618 149546 115174
rect 150102 114618 185546 115174
rect 186102 114618 221546 115174
rect 222102 114618 257546 115174
rect 258102 114618 293546 115174
rect 294102 114618 329546 115174
rect 330102 114618 365546 115174
rect 366102 114618 401546 115174
rect 402102 114618 437546 115174
rect 438102 114618 473546 115174
rect 474102 114618 509546 115174
rect 510102 114618 545546 115174
rect 546102 114618 581546 115174
rect 582102 114618 587262 115174
rect 587818 114618 588810 115174
rect -4886 114586 588810 114618
rect -2966 111454 586890 111486
rect -2966 110898 -1974 111454
rect -1418 110898 1826 111454
rect 2382 110898 37826 111454
rect 38382 110898 73826 111454
rect 74382 110898 109826 111454
rect 110382 110898 145826 111454
rect 146382 110898 181826 111454
rect 182382 110898 217826 111454
rect 218382 110898 253826 111454
rect 254382 110898 289826 111454
rect 290382 110898 325826 111454
rect 326382 110898 361826 111454
rect 362382 110898 397826 111454
rect 398382 110898 433826 111454
rect 434382 110898 469826 111454
rect 470382 110898 505826 111454
rect 506382 110898 541826 111454
rect 542382 110898 577826 111454
rect 578382 110898 585342 111454
rect 585898 110898 586890 111454
rect -2966 110866 586890 110898
rect -8726 104614 592650 104646
rect -8726 104058 -8694 104614
rect -8138 104058 30986 104614
rect 31542 104058 66986 104614
rect 67542 104058 102986 104614
rect 103542 104058 138986 104614
rect 139542 104058 174986 104614
rect 175542 104058 210986 104614
rect 211542 104058 246986 104614
rect 247542 104058 282986 104614
rect 283542 104058 318986 104614
rect 319542 104058 354986 104614
rect 355542 104058 390986 104614
rect 391542 104058 426986 104614
rect 427542 104058 462986 104614
rect 463542 104058 498986 104614
rect 499542 104058 534986 104614
rect 535542 104058 570986 104614
rect 571542 104058 592062 104614
rect 592618 104058 592650 104614
rect -8726 104026 592650 104058
rect -6806 100894 590730 100926
rect -6806 100338 -6774 100894
rect -6218 100338 27266 100894
rect 27822 100338 63266 100894
rect 63822 100338 99266 100894
rect 99822 100338 135266 100894
rect 135822 100338 171266 100894
rect 171822 100338 207266 100894
rect 207822 100338 243266 100894
rect 243822 100338 279266 100894
rect 279822 100338 315266 100894
rect 315822 100338 351266 100894
rect 351822 100338 387266 100894
rect 387822 100338 423266 100894
rect 423822 100338 459266 100894
rect 459822 100338 495266 100894
rect 495822 100338 531266 100894
rect 531822 100338 567266 100894
rect 567822 100338 590142 100894
rect 590698 100338 590730 100894
rect -6806 100306 590730 100338
rect -4886 97174 588810 97206
rect -4886 96618 -4854 97174
rect -4298 96618 23546 97174
rect 24102 96618 59546 97174
rect 60102 96618 95546 97174
rect 96102 96618 131546 97174
rect 132102 96618 167546 97174
rect 168102 96618 203546 97174
rect 204102 96618 239546 97174
rect 240102 96618 275546 97174
rect 276102 96618 311546 97174
rect 312102 96618 347546 97174
rect 348102 96618 383546 97174
rect 384102 96618 419546 97174
rect 420102 96618 455546 97174
rect 456102 96618 491546 97174
rect 492102 96618 527546 97174
rect 528102 96618 563546 97174
rect 564102 96618 588222 97174
rect 588778 96618 588810 97174
rect -4886 96586 588810 96618
rect -2966 93454 586890 93486
rect -2966 92898 -2934 93454
rect -2378 92898 19826 93454
rect 20382 92898 55826 93454
rect 56382 92898 91826 93454
rect 92382 92898 127826 93454
rect 128382 92898 163826 93454
rect 164382 92898 199826 93454
rect 200382 92898 235826 93454
rect 236382 92898 271826 93454
rect 272382 92898 307826 93454
rect 308382 92898 343826 93454
rect 344382 92898 379826 93454
rect 380382 92898 415826 93454
rect 416382 92898 451826 93454
rect 452382 92898 487826 93454
rect 488382 92898 523826 93454
rect 524382 92898 559826 93454
rect 560382 92898 586302 93454
rect 586858 92898 586890 93454
rect -2966 92866 586890 92898
rect -8726 86614 592650 86646
rect -8726 86058 -7734 86614
rect -7178 86058 12986 86614
rect 13542 86058 48986 86614
rect 49542 86058 84986 86614
rect 85542 86058 120986 86614
rect 121542 86058 156986 86614
rect 157542 86058 192986 86614
rect 193542 86058 228986 86614
rect 229542 86058 264986 86614
rect 265542 86058 300986 86614
rect 301542 86058 336986 86614
rect 337542 86058 372986 86614
rect 373542 86058 408986 86614
rect 409542 86058 444986 86614
rect 445542 86058 480986 86614
rect 481542 86058 516986 86614
rect 517542 86058 552986 86614
rect 553542 86058 591102 86614
rect 591658 86058 592650 86614
rect -8726 86026 592650 86058
rect -6806 82894 590730 82926
rect -6806 82338 -5814 82894
rect -5258 82338 9266 82894
rect 9822 82338 45266 82894
rect 45822 82338 81266 82894
rect 81822 82338 117266 82894
rect 117822 82338 153266 82894
rect 153822 82338 189266 82894
rect 189822 82338 225266 82894
rect 225822 82338 261266 82894
rect 261822 82338 297266 82894
rect 297822 82338 333266 82894
rect 333822 82338 369266 82894
rect 369822 82338 405266 82894
rect 405822 82338 441266 82894
rect 441822 82338 477266 82894
rect 477822 82338 513266 82894
rect 513822 82338 549266 82894
rect 549822 82338 589182 82894
rect 589738 82338 590730 82894
rect -6806 82306 590730 82338
rect -4886 79174 588810 79206
rect -4886 78618 -3894 79174
rect -3338 78618 5546 79174
rect 6102 78618 41546 79174
rect 42102 78618 77546 79174
rect 78102 78618 113546 79174
rect 114102 78618 149546 79174
rect 150102 78618 185546 79174
rect 186102 78618 221546 79174
rect 222102 78618 257546 79174
rect 258102 78618 293546 79174
rect 294102 78618 329546 79174
rect 330102 78618 365546 79174
rect 366102 78618 401546 79174
rect 402102 78618 437546 79174
rect 438102 78618 473546 79174
rect 474102 78618 509546 79174
rect 510102 78618 545546 79174
rect 546102 78618 581546 79174
rect 582102 78618 587262 79174
rect 587818 78618 588810 79174
rect -4886 78586 588810 78618
rect -2966 75454 586890 75486
rect -2966 74898 -1974 75454
rect -1418 74898 1826 75454
rect 2382 74898 37826 75454
rect 38382 74898 73826 75454
rect 74382 74898 109826 75454
rect 110382 74898 145826 75454
rect 146382 74898 181826 75454
rect 182382 74898 217826 75454
rect 218382 74898 253826 75454
rect 254382 74898 289826 75454
rect 290382 74898 325826 75454
rect 326382 74898 361826 75454
rect 362382 74898 397826 75454
rect 398382 74898 433826 75454
rect 434382 74898 469826 75454
rect 470382 74898 505826 75454
rect 506382 74898 541826 75454
rect 542382 74898 577826 75454
rect 578382 74898 585342 75454
rect 585898 74898 586890 75454
rect -2966 74866 586890 74898
rect -8726 68614 592650 68646
rect -8726 68058 -8694 68614
rect -8138 68058 30986 68614
rect 31542 68058 66986 68614
rect 67542 68058 102986 68614
rect 103542 68058 138986 68614
rect 139542 68058 174986 68614
rect 175542 68058 210986 68614
rect 211542 68058 246986 68614
rect 247542 68058 282986 68614
rect 283542 68058 318986 68614
rect 319542 68058 354986 68614
rect 355542 68058 390986 68614
rect 391542 68058 426986 68614
rect 427542 68058 462986 68614
rect 463542 68058 498986 68614
rect 499542 68058 534986 68614
rect 535542 68058 570986 68614
rect 571542 68058 592062 68614
rect 592618 68058 592650 68614
rect -8726 68026 592650 68058
rect -6806 64894 590730 64926
rect -6806 64338 -6774 64894
rect -6218 64338 27266 64894
rect 27822 64338 63266 64894
rect 63822 64338 99266 64894
rect 99822 64338 135266 64894
rect 135822 64338 171266 64894
rect 171822 64338 207266 64894
rect 207822 64338 243266 64894
rect 243822 64338 279266 64894
rect 279822 64338 315266 64894
rect 315822 64338 351266 64894
rect 351822 64338 387266 64894
rect 387822 64338 423266 64894
rect 423822 64338 459266 64894
rect 459822 64338 495266 64894
rect 495822 64338 531266 64894
rect 531822 64338 567266 64894
rect 567822 64338 590142 64894
rect 590698 64338 590730 64894
rect -6806 64306 590730 64338
rect -4886 61174 588810 61206
rect -4886 60618 -4854 61174
rect -4298 60618 23546 61174
rect 24102 60618 59546 61174
rect 60102 60618 95546 61174
rect 96102 60618 131546 61174
rect 132102 60618 167546 61174
rect 168102 60618 203546 61174
rect 204102 60618 239546 61174
rect 240102 60618 275546 61174
rect 276102 60618 311546 61174
rect 312102 60618 347546 61174
rect 348102 60618 383546 61174
rect 384102 60618 419546 61174
rect 420102 60618 455546 61174
rect 456102 60618 491546 61174
rect 492102 60618 527546 61174
rect 528102 60618 563546 61174
rect 564102 60618 588222 61174
rect 588778 60618 588810 61174
rect -4886 60586 588810 60618
rect -2966 57454 586890 57486
rect -2966 56898 -2934 57454
rect -2378 56898 19826 57454
rect 20382 56898 55826 57454
rect 56382 56898 91826 57454
rect 92382 56898 127826 57454
rect 128382 56898 163826 57454
rect 164382 56898 199826 57454
rect 200382 56898 235826 57454
rect 236382 56898 271826 57454
rect 272382 56898 307826 57454
rect 308382 56898 343826 57454
rect 344382 56898 379826 57454
rect 380382 56898 415826 57454
rect 416382 56898 451826 57454
rect 452382 56898 487826 57454
rect 488382 56898 523826 57454
rect 524382 56898 559826 57454
rect 560382 56898 586302 57454
rect 586858 56898 586890 57454
rect -2966 56866 586890 56898
rect -8726 50614 592650 50646
rect -8726 50058 -7734 50614
rect -7178 50058 12986 50614
rect 13542 50058 48986 50614
rect 49542 50058 84986 50614
rect 85542 50058 120986 50614
rect 121542 50058 156986 50614
rect 157542 50058 192986 50614
rect 193542 50058 228986 50614
rect 229542 50058 264986 50614
rect 265542 50058 300986 50614
rect 301542 50058 336986 50614
rect 337542 50058 372986 50614
rect 373542 50058 408986 50614
rect 409542 50058 444986 50614
rect 445542 50058 480986 50614
rect 481542 50058 516986 50614
rect 517542 50058 552986 50614
rect 553542 50058 591102 50614
rect 591658 50058 592650 50614
rect -8726 50026 592650 50058
rect -6806 46894 590730 46926
rect -6806 46338 -5814 46894
rect -5258 46338 9266 46894
rect 9822 46338 45266 46894
rect 45822 46338 81266 46894
rect 81822 46338 117266 46894
rect 117822 46338 153266 46894
rect 153822 46338 189266 46894
rect 189822 46338 225266 46894
rect 225822 46338 261266 46894
rect 261822 46338 297266 46894
rect 297822 46338 333266 46894
rect 333822 46338 369266 46894
rect 369822 46338 405266 46894
rect 405822 46338 441266 46894
rect 441822 46338 477266 46894
rect 477822 46338 513266 46894
rect 513822 46338 549266 46894
rect 549822 46338 589182 46894
rect 589738 46338 590730 46894
rect -6806 46306 590730 46338
rect -4886 43174 588810 43206
rect -4886 42618 -3894 43174
rect -3338 42618 5546 43174
rect 6102 42618 41546 43174
rect 42102 42618 77546 43174
rect 78102 42618 113546 43174
rect 114102 42618 149546 43174
rect 150102 42618 185546 43174
rect 186102 42618 221546 43174
rect 222102 42618 257546 43174
rect 258102 42618 293546 43174
rect 294102 42618 329546 43174
rect 330102 42618 365546 43174
rect 366102 42618 401546 43174
rect 402102 42618 437546 43174
rect 438102 42618 473546 43174
rect 474102 42618 509546 43174
rect 510102 42618 545546 43174
rect 546102 42618 581546 43174
rect 582102 42618 587262 43174
rect 587818 42618 588810 43174
rect -4886 42586 588810 42618
rect -2966 39454 586890 39486
rect -2966 38898 -1974 39454
rect -1418 38898 1826 39454
rect 2382 38898 37826 39454
rect 38382 38898 73826 39454
rect 74382 38898 109826 39454
rect 110382 38898 145826 39454
rect 146382 38898 181826 39454
rect 182382 38898 217826 39454
rect 218382 38898 253826 39454
rect 254382 38898 289826 39454
rect 290382 38898 325826 39454
rect 326382 38898 361826 39454
rect 362382 38898 397826 39454
rect 398382 38898 433826 39454
rect 434382 38898 469826 39454
rect 470382 38898 505826 39454
rect 506382 38898 541826 39454
rect 542382 38898 577826 39454
rect 578382 38898 585342 39454
rect 585898 38898 586890 39454
rect -2966 38866 586890 38898
rect -8726 32614 592650 32646
rect -8726 32058 -8694 32614
rect -8138 32058 30986 32614
rect 31542 32058 66986 32614
rect 67542 32058 102986 32614
rect 103542 32058 138986 32614
rect 139542 32058 174986 32614
rect 175542 32058 210986 32614
rect 211542 32058 246986 32614
rect 247542 32058 282986 32614
rect 283542 32058 318986 32614
rect 319542 32058 354986 32614
rect 355542 32058 390986 32614
rect 391542 32058 426986 32614
rect 427542 32058 462986 32614
rect 463542 32058 498986 32614
rect 499542 32058 534986 32614
rect 535542 32058 570986 32614
rect 571542 32058 592062 32614
rect 592618 32058 592650 32614
rect -8726 32026 592650 32058
rect -6806 28894 590730 28926
rect -6806 28338 -6774 28894
rect -6218 28338 27266 28894
rect 27822 28338 63266 28894
rect 63822 28338 99266 28894
rect 99822 28338 135266 28894
rect 135822 28338 171266 28894
rect 171822 28338 207266 28894
rect 207822 28338 243266 28894
rect 243822 28338 279266 28894
rect 279822 28338 315266 28894
rect 315822 28338 351266 28894
rect 351822 28338 387266 28894
rect 387822 28338 423266 28894
rect 423822 28338 459266 28894
rect 459822 28338 495266 28894
rect 495822 28338 531266 28894
rect 531822 28338 567266 28894
rect 567822 28338 590142 28894
rect 590698 28338 590730 28894
rect -6806 28306 590730 28338
rect -4886 25174 588810 25206
rect -4886 24618 -4854 25174
rect -4298 24618 23546 25174
rect 24102 24618 59546 25174
rect 60102 24618 95546 25174
rect 96102 24618 131546 25174
rect 132102 24618 167546 25174
rect 168102 24618 203546 25174
rect 204102 24618 239546 25174
rect 240102 24618 275546 25174
rect 276102 24618 311546 25174
rect 312102 24618 347546 25174
rect 348102 24618 383546 25174
rect 384102 24618 419546 25174
rect 420102 24618 455546 25174
rect 456102 24618 491546 25174
rect 492102 24618 527546 25174
rect 528102 24618 563546 25174
rect 564102 24618 588222 25174
rect 588778 24618 588810 25174
rect -4886 24586 588810 24618
rect -2966 21454 586890 21486
rect -2966 20898 -2934 21454
rect -2378 20898 19826 21454
rect 20382 20898 55826 21454
rect 56382 20898 91826 21454
rect 92382 20898 127826 21454
rect 128382 20898 163826 21454
rect 164382 20898 199826 21454
rect 200382 20898 235826 21454
rect 236382 20898 271826 21454
rect 272382 20898 307826 21454
rect 308382 20898 343826 21454
rect 344382 20898 379826 21454
rect 380382 20898 415826 21454
rect 416382 20898 451826 21454
rect 452382 20898 487826 21454
rect 488382 20898 523826 21454
rect 524382 20898 559826 21454
rect 560382 20898 586302 21454
rect 586858 20898 586890 21454
rect -2966 20866 586890 20898
rect -8726 14614 592650 14646
rect -8726 14058 -7734 14614
rect -7178 14058 12986 14614
rect 13542 14058 48986 14614
rect 49542 14058 84986 14614
rect 85542 14058 120986 14614
rect 121542 14058 156986 14614
rect 157542 14058 192986 14614
rect 193542 14058 228986 14614
rect 229542 14058 264986 14614
rect 265542 14058 300986 14614
rect 301542 14058 336986 14614
rect 337542 14058 372986 14614
rect 373542 14058 408986 14614
rect 409542 14058 444986 14614
rect 445542 14058 480986 14614
rect 481542 14058 516986 14614
rect 517542 14058 552986 14614
rect 553542 14058 591102 14614
rect 591658 14058 592650 14614
rect -8726 14026 592650 14058
rect -6806 10894 590730 10926
rect -6806 10338 -5814 10894
rect -5258 10338 9266 10894
rect 9822 10338 45266 10894
rect 45822 10338 81266 10894
rect 81822 10338 117266 10894
rect 117822 10338 153266 10894
rect 153822 10338 189266 10894
rect 189822 10338 225266 10894
rect 225822 10338 261266 10894
rect 261822 10338 297266 10894
rect 297822 10338 333266 10894
rect 333822 10338 369266 10894
rect 369822 10338 405266 10894
rect 405822 10338 441266 10894
rect 441822 10338 477266 10894
rect 477822 10338 513266 10894
rect 513822 10338 549266 10894
rect 549822 10338 589182 10894
rect 589738 10338 590730 10894
rect -6806 10306 590730 10338
rect -4886 7174 588810 7206
rect -4886 6618 -3894 7174
rect -3338 6618 5546 7174
rect 6102 6618 41546 7174
rect 42102 6618 77546 7174
rect 78102 6618 113546 7174
rect 114102 6618 149546 7174
rect 150102 6618 185546 7174
rect 186102 6618 221546 7174
rect 222102 6618 257546 7174
rect 258102 6618 293546 7174
rect 294102 6618 329546 7174
rect 330102 6618 365546 7174
rect 366102 6618 401546 7174
rect 402102 6618 437546 7174
rect 438102 6618 473546 7174
rect 474102 6618 509546 7174
rect 510102 6618 545546 7174
rect 546102 6618 581546 7174
rect 582102 6618 587262 7174
rect 587818 6618 588810 7174
rect -4886 6586 588810 6618
rect -2966 3454 586890 3486
rect -2966 2898 -1974 3454
rect -1418 2898 1826 3454
rect 2382 2898 37826 3454
rect 38382 2898 73826 3454
rect 74382 2898 109826 3454
rect 110382 2898 145826 3454
rect 146382 2898 181826 3454
rect 182382 2898 217826 3454
rect 218382 2898 253826 3454
rect 254382 2898 289826 3454
rect 290382 2898 325826 3454
rect 326382 2898 361826 3454
rect 362382 2898 397826 3454
rect 398382 2898 433826 3454
rect 434382 2898 469826 3454
rect 470382 2898 505826 3454
rect 506382 2898 541826 3454
rect 542382 2898 577826 3454
rect 578382 2898 585342 3454
rect 585898 2898 586890 3454
rect -2966 2866 586890 2898
rect -2006 -346 585930 -314
rect -2006 -902 -1974 -346
rect -1418 -902 1826 -346
rect 2382 -902 37826 -346
rect 38382 -902 73826 -346
rect 74382 -902 109826 -346
rect 110382 -902 145826 -346
rect 146382 -902 181826 -346
rect 182382 -902 217826 -346
rect 218382 -902 253826 -346
rect 254382 -902 289826 -346
rect 290382 -902 325826 -346
rect 326382 -902 361826 -346
rect 362382 -902 397826 -346
rect 398382 -902 433826 -346
rect 434382 -902 469826 -346
rect 470382 -902 505826 -346
rect 506382 -902 541826 -346
rect 542382 -902 577826 -346
rect 578382 -902 585342 -346
rect 585898 -902 585930 -346
rect -2006 -934 585930 -902
rect -2966 -1306 586890 -1274
rect -2966 -1862 -2934 -1306
rect -2378 -1862 19826 -1306
rect 20382 -1862 55826 -1306
rect 56382 -1862 91826 -1306
rect 92382 -1862 127826 -1306
rect 128382 -1862 163826 -1306
rect 164382 -1862 199826 -1306
rect 200382 -1862 235826 -1306
rect 236382 -1862 271826 -1306
rect 272382 -1862 307826 -1306
rect 308382 -1862 343826 -1306
rect 344382 -1862 379826 -1306
rect 380382 -1862 415826 -1306
rect 416382 -1862 451826 -1306
rect 452382 -1862 487826 -1306
rect 488382 -1862 523826 -1306
rect 524382 -1862 559826 -1306
rect 560382 -1862 586302 -1306
rect 586858 -1862 586890 -1306
rect -2966 -1894 586890 -1862
rect -3926 -2266 587850 -2234
rect -3926 -2822 -3894 -2266
rect -3338 -2822 5546 -2266
rect 6102 -2822 41546 -2266
rect 42102 -2822 77546 -2266
rect 78102 -2822 113546 -2266
rect 114102 -2822 149546 -2266
rect 150102 -2822 185546 -2266
rect 186102 -2822 221546 -2266
rect 222102 -2822 257546 -2266
rect 258102 -2822 293546 -2266
rect 294102 -2822 329546 -2266
rect 330102 -2822 365546 -2266
rect 366102 -2822 401546 -2266
rect 402102 -2822 437546 -2266
rect 438102 -2822 473546 -2266
rect 474102 -2822 509546 -2266
rect 510102 -2822 545546 -2266
rect 546102 -2822 581546 -2266
rect 582102 -2822 587262 -2266
rect 587818 -2822 587850 -2266
rect -3926 -2854 587850 -2822
rect -4886 -3226 588810 -3194
rect -4886 -3782 -4854 -3226
rect -4298 -3782 23546 -3226
rect 24102 -3782 59546 -3226
rect 60102 -3782 95546 -3226
rect 96102 -3782 131546 -3226
rect 132102 -3782 167546 -3226
rect 168102 -3782 203546 -3226
rect 204102 -3782 239546 -3226
rect 240102 -3782 275546 -3226
rect 276102 -3782 311546 -3226
rect 312102 -3782 347546 -3226
rect 348102 -3782 383546 -3226
rect 384102 -3782 419546 -3226
rect 420102 -3782 455546 -3226
rect 456102 -3782 491546 -3226
rect 492102 -3782 527546 -3226
rect 528102 -3782 563546 -3226
rect 564102 -3782 588222 -3226
rect 588778 -3782 588810 -3226
rect -4886 -3814 588810 -3782
rect -5846 -4186 589770 -4154
rect -5846 -4742 -5814 -4186
rect -5258 -4742 9266 -4186
rect 9822 -4742 45266 -4186
rect 45822 -4742 81266 -4186
rect 81822 -4742 117266 -4186
rect 117822 -4742 153266 -4186
rect 153822 -4742 189266 -4186
rect 189822 -4742 225266 -4186
rect 225822 -4742 261266 -4186
rect 261822 -4742 297266 -4186
rect 297822 -4742 333266 -4186
rect 333822 -4742 369266 -4186
rect 369822 -4742 405266 -4186
rect 405822 -4742 441266 -4186
rect 441822 -4742 477266 -4186
rect 477822 -4742 513266 -4186
rect 513822 -4742 549266 -4186
rect 549822 -4742 589182 -4186
rect 589738 -4742 589770 -4186
rect -5846 -4774 589770 -4742
rect -6806 -5146 590730 -5114
rect -6806 -5702 -6774 -5146
rect -6218 -5702 27266 -5146
rect 27822 -5702 63266 -5146
rect 63822 -5702 99266 -5146
rect 99822 -5702 135266 -5146
rect 135822 -5702 171266 -5146
rect 171822 -5702 207266 -5146
rect 207822 -5702 243266 -5146
rect 243822 -5702 279266 -5146
rect 279822 -5702 315266 -5146
rect 315822 -5702 351266 -5146
rect 351822 -5702 387266 -5146
rect 387822 -5702 423266 -5146
rect 423822 -5702 459266 -5146
rect 459822 -5702 495266 -5146
rect 495822 -5702 531266 -5146
rect 531822 -5702 567266 -5146
rect 567822 -5702 590142 -5146
rect 590698 -5702 590730 -5146
rect -6806 -5734 590730 -5702
rect -7766 -6106 591690 -6074
rect -7766 -6662 -7734 -6106
rect -7178 -6662 12986 -6106
rect 13542 -6662 48986 -6106
rect 49542 -6662 84986 -6106
rect 85542 -6662 120986 -6106
rect 121542 -6662 156986 -6106
rect 157542 -6662 192986 -6106
rect 193542 -6662 228986 -6106
rect 229542 -6662 264986 -6106
rect 265542 -6662 300986 -6106
rect 301542 -6662 336986 -6106
rect 337542 -6662 372986 -6106
rect 373542 -6662 408986 -6106
rect 409542 -6662 444986 -6106
rect 445542 -6662 480986 -6106
rect 481542 -6662 516986 -6106
rect 517542 -6662 552986 -6106
rect 553542 -6662 591102 -6106
rect 591658 -6662 591690 -6106
rect -7766 -6694 591690 -6662
rect -8726 -7066 592650 -7034
rect -8726 -7622 -8694 -7066
rect -8138 -7622 30986 -7066
rect 31542 -7622 66986 -7066
rect 67542 -7622 102986 -7066
rect 103542 -7622 138986 -7066
rect 139542 -7622 174986 -7066
rect 175542 -7622 210986 -7066
rect 211542 -7622 246986 -7066
rect 247542 -7622 282986 -7066
rect 283542 -7622 318986 -7066
rect 319542 -7622 354986 -7066
rect 355542 -7622 390986 -7066
rect 391542 -7622 426986 -7066
rect 427542 -7622 462986 -7066
rect 463542 -7622 498986 -7066
rect 499542 -7622 534986 -7066
rect 535542 -7622 570986 -7066
rect 571542 -7622 592062 -7066
rect 592618 -7622 592650 -7066
rect -8726 -7654 592650 -7622
use user_proj_example  mprj
timestamp 1639277212
transform 1 0 235000 0 1 338000
box 106 0 147278 149603
<< labels >>
rlabel metal3 s 583520 285276 584960 285516 4 analog_io[0]
port 1 nsew
rlabel metal2 s 446098 703520 446210 704960 4 analog_io[10]
port 2 nsew
rlabel metal2 s 381146 703520 381258 704960 4 analog_io[11]
port 3 nsew
rlabel metal2 s 316286 703520 316398 704960 4 analog_io[12]
port 4 nsew
rlabel metal2 s 251426 703520 251538 704960 4 analog_io[13]
port 5 nsew
rlabel metal2 s 186474 703520 186586 704960 4 analog_io[14]
port 6 nsew
rlabel metal2 s 121614 703520 121726 704960 4 analog_io[15]
port 7 nsew
rlabel metal2 s 56754 703520 56866 704960 4 analog_io[16]
port 8 nsew
rlabel metal3 s -960 697220 480 697460 4 analog_io[17]
port 9 nsew
rlabel metal3 s -960 644996 480 645236 4 analog_io[18]
port 10 nsew
rlabel metal3 s -960 592908 480 593148 4 analog_io[19]
port 11 nsew
rlabel metal3 s 583520 338452 584960 338692 4 analog_io[1]
port 12 nsew
rlabel metal3 s -960 540684 480 540924 4 analog_io[20]
port 13 nsew
rlabel metal3 s -960 488596 480 488836 4 analog_io[21]
port 14 nsew
rlabel metal3 s -960 436508 480 436748 4 analog_io[22]
port 15 nsew
rlabel metal3 s -960 384284 480 384524 4 analog_io[23]
port 16 nsew
rlabel metal3 s -960 332196 480 332436 4 analog_io[24]
port 17 nsew
rlabel metal3 s -960 279972 480 280212 4 analog_io[25]
port 18 nsew
rlabel metal3 s -960 227884 480 228124 4 analog_io[26]
port 19 nsew
rlabel metal3 s -960 175796 480 176036 4 analog_io[27]
port 20 nsew
rlabel metal3 s -960 123572 480 123812 4 analog_io[28]
port 21 nsew
rlabel metal3 s 583520 391628 584960 391868 4 analog_io[2]
port 22 nsew
rlabel metal3 s 583520 444668 584960 444908 4 analog_io[3]
port 23 nsew
rlabel metal3 s 583520 497844 584960 498084 4 analog_io[4]
port 24 nsew
rlabel metal3 s 583520 551020 584960 551260 4 analog_io[5]
port 25 nsew
rlabel metal3 s 583520 604060 584960 604300 4 analog_io[6]
port 26 nsew
rlabel metal3 s 583520 657236 584960 657476 4 analog_io[7]
port 27 nsew
rlabel metal2 s 575818 703520 575930 704960 4 analog_io[8]
port 28 nsew
rlabel metal2 s 510958 703520 511070 704960 4 analog_io[9]
port 29 nsew
rlabel metal3 s 583520 6476 584960 6716 4 io_in[0]
port 30 nsew
rlabel metal3 s 583520 457996 584960 458236 4 io_in[10]
port 31 nsew
rlabel metal3 s 583520 511172 584960 511412 4 io_in[11]
port 32 nsew
rlabel metal3 s 583520 564212 584960 564452 4 io_in[12]
port 33 nsew
rlabel metal3 s 583520 617388 584960 617628 4 io_in[13]
port 34 nsew
rlabel metal3 s 583520 670564 584960 670804 4 io_in[14]
port 35 nsew
rlabel metal2 s 559626 703520 559738 704960 4 io_in[15]
port 36 nsew
rlabel metal2 s 494766 703520 494878 704960 4 io_in[16]
port 37 nsew
rlabel metal2 s 429814 703520 429926 704960 4 io_in[17]
port 38 nsew
rlabel metal2 s 364954 703520 365066 704960 4 io_in[18]
port 39 nsew
rlabel metal2 s 300094 703520 300206 704960 4 io_in[19]
port 40 nsew
rlabel metal3 s 583520 46188 584960 46428 4 io_in[1]
port 41 nsew
rlabel metal2 s 235142 703520 235254 704960 4 io_in[20]
port 42 nsew
rlabel metal2 s 170282 703520 170394 704960 4 io_in[21]
port 43 nsew
rlabel metal2 s 105422 703520 105534 704960 4 io_in[22]
port 44 nsew
rlabel metal2 s 40470 703520 40582 704960 4 io_in[23]
port 45 nsew
rlabel metal3 s -960 684164 480 684404 4 io_in[24]
port 46 nsew
rlabel metal3 s -960 631940 480 632180 4 io_in[25]
port 47 nsew
rlabel metal3 s -960 579852 480 580092 4 io_in[26]
port 48 nsew
rlabel metal3 s -960 527764 480 528004 4 io_in[27]
port 49 nsew
rlabel metal3 s -960 475540 480 475780 4 io_in[28]
port 50 nsew
rlabel metal3 s -960 423452 480 423692 4 io_in[29]
port 51 nsew
rlabel metal3 s 583520 86036 584960 86276 4 io_in[2]
port 52 nsew
rlabel metal3 s -960 371228 480 371468 4 io_in[30]
port 53 nsew
rlabel metal3 s -960 319140 480 319380 4 io_in[31]
port 54 nsew
rlabel metal3 s -960 267052 480 267292 4 io_in[32]
port 55 nsew
rlabel metal3 s -960 214828 480 215068 4 io_in[33]
port 56 nsew
rlabel metal3 s -960 162740 480 162980 4 io_in[34]
port 57 nsew
rlabel metal3 s -960 110516 480 110756 4 io_in[35]
port 58 nsew
rlabel metal3 s -960 71484 480 71724 4 io_in[36]
port 59 nsew
rlabel metal3 s -960 32316 480 32556 4 io_in[37]
port 60 nsew
rlabel metal3 s 583520 125884 584960 126124 4 io_in[3]
port 61 nsew
rlabel metal3 s 583520 165732 584960 165972 4 io_in[4]
port 62 nsew
rlabel metal3 s 583520 205580 584960 205820 4 io_in[5]
port 63 nsew
rlabel metal3 s 583520 245428 584960 245668 4 io_in[6]
port 64 nsew
rlabel metal3 s 583520 298604 584960 298844 4 io_in[7]
port 65 nsew
rlabel metal3 s 583520 351780 584960 352020 4 io_in[8]
port 66 nsew
rlabel metal3 s 583520 404820 584960 405060 4 io_in[9]
port 67 nsew
rlabel metal3 s 583520 32996 584960 33236 4 io_oeb[0]
port 68 nsew
rlabel metal3 s 583520 484516 584960 484756 4 io_oeb[10]
port 69 nsew
rlabel metal3 s 583520 537692 584960 537932 4 io_oeb[11]
port 70 nsew
rlabel metal3 s 583520 590868 584960 591108 4 io_oeb[12]
port 71 nsew
rlabel metal3 s 583520 643908 584960 644148 4 io_oeb[13]
port 72 nsew
rlabel metal3 s 583520 697084 584960 697324 4 io_oeb[14]
port 73 nsew
rlabel metal2 s 527150 703520 527262 704960 4 io_oeb[15]
port 74 nsew
rlabel metal2 s 462290 703520 462402 704960 4 io_oeb[16]
port 75 nsew
rlabel metal2 s 397430 703520 397542 704960 4 io_oeb[17]
port 76 nsew
rlabel metal2 s 332478 703520 332590 704960 4 io_oeb[18]
port 77 nsew
rlabel metal2 s 267618 703520 267730 704960 4 io_oeb[19]
port 78 nsew
rlabel metal3 s 583520 72844 584960 73084 4 io_oeb[1]
port 79 nsew
rlabel metal2 s 202758 703520 202870 704960 4 io_oeb[20]
port 80 nsew
rlabel metal2 s 137806 703520 137918 704960 4 io_oeb[21]
port 81 nsew
rlabel metal2 s 72946 703520 73058 704960 4 io_oeb[22]
port 82 nsew
rlabel metal2 s 8086 703520 8198 704960 4 io_oeb[23]
port 83 nsew
rlabel metal3 s -960 658052 480 658292 4 io_oeb[24]
port 84 nsew
rlabel metal3 s -960 605964 480 606204 4 io_oeb[25]
port 85 nsew
rlabel metal3 s -960 553740 480 553980 4 io_oeb[26]
port 86 nsew
rlabel metal3 s -960 501652 480 501892 4 io_oeb[27]
port 87 nsew
rlabel metal3 s -960 449428 480 449668 4 io_oeb[28]
port 88 nsew
rlabel metal3 s -960 397340 480 397580 4 io_oeb[29]
port 89 nsew
rlabel metal3 s 583520 112692 584960 112932 4 io_oeb[2]
port 90 nsew
rlabel metal3 s -960 345252 480 345492 4 io_oeb[30]
port 91 nsew
rlabel metal3 s -960 293028 480 293268 4 io_oeb[31]
port 92 nsew
rlabel metal3 s -960 240940 480 241180 4 io_oeb[32]
port 93 nsew
rlabel metal3 s -960 188716 480 188956 4 io_oeb[33]
port 94 nsew
rlabel metal3 s -960 136628 480 136868 4 io_oeb[34]
port 95 nsew
rlabel metal3 s -960 84540 480 84780 4 io_oeb[35]
port 96 nsew
rlabel metal3 s -960 45372 480 45612 4 io_oeb[36]
port 97 nsew
rlabel metal3 s -960 6340 480 6580 4 io_oeb[37]
port 98 nsew
rlabel metal3 s 583520 152540 584960 152780 4 io_oeb[3]
port 99 nsew
rlabel metal3 s 583520 192388 584960 192628 4 io_oeb[4]
port 100 nsew
rlabel metal3 s 583520 232236 584960 232476 4 io_oeb[5]
port 101 nsew
rlabel metal3 s 583520 272084 584960 272324 4 io_oeb[6]
port 102 nsew
rlabel metal3 s 583520 325124 584960 325364 4 io_oeb[7]
port 103 nsew
rlabel metal3 s 583520 378300 584960 378540 4 io_oeb[8]
port 104 nsew
rlabel metal3 s 583520 431476 584960 431716 4 io_oeb[9]
port 105 nsew
rlabel metal3 s 583520 19668 584960 19908 4 io_out[0]
port 106 nsew
rlabel metal3 s 583520 471324 584960 471564 4 io_out[10]
port 107 nsew
rlabel metal3 s 583520 524364 584960 524604 4 io_out[11]
port 108 nsew
rlabel metal3 s 583520 577540 584960 577780 4 io_out[12]
port 109 nsew
rlabel metal3 s 583520 630716 584960 630956 4 io_out[13]
port 110 nsew
rlabel metal3 s 583520 683756 584960 683996 4 io_out[14]
port 111 nsew
rlabel metal2 s 543434 703520 543546 704960 4 io_out[15]
port 112 nsew
rlabel metal2 s 478482 703520 478594 704960 4 io_out[16]
port 113 nsew
rlabel metal2 s 413622 703520 413734 704960 4 io_out[17]
port 114 nsew
rlabel metal2 s 348762 703520 348874 704960 4 io_out[18]
port 115 nsew
rlabel metal2 s 283810 703520 283922 704960 4 io_out[19]
port 116 nsew
rlabel metal3 s 583520 59516 584960 59756 4 io_out[1]
port 117 nsew
rlabel metal2 s 218950 703520 219062 704960 4 io_out[20]
port 118 nsew
rlabel metal2 s 154090 703520 154202 704960 4 io_out[21]
port 119 nsew
rlabel metal2 s 89138 703520 89250 704960 4 io_out[22]
port 120 nsew
rlabel metal2 s 24278 703520 24390 704960 4 io_out[23]
port 121 nsew
rlabel metal3 s -960 671108 480 671348 4 io_out[24]
port 122 nsew
rlabel metal3 s -960 619020 480 619260 4 io_out[25]
port 123 nsew
rlabel metal3 s -960 566796 480 567036 4 io_out[26]
port 124 nsew
rlabel metal3 s -960 514708 480 514948 4 io_out[27]
port 125 nsew
rlabel metal3 s -960 462484 480 462724 4 io_out[28]
port 126 nsew
rlabel metal3 s -960 410396 480 410636 4 io_out[29]
port 127 nsew
rlabel metal3 s 583520 99364 584960 99604 4 io_out[2]
port 128 nsew
rlabel metal3 s -960 358308 480 358548 4 io_out[30]
port 129 nsew
rlabel metal3 s -960 306084 480 306324 4 io_out[31]
port 130 nsew
rlabel metal3 s -960 253996 480 254236 4 io_out[32]
port 131 nsew
rlabel metal3 s -960 201772 480 202012 4 io_out[33]
port 132 nsew
rlabel metal3 s -960 149684 480 149924 4 io_out[34]
port 133 nsew
rlabel metal3 s -960 97460 480 97700 4 io_out[35]
port 134 nsew
rlabel metal3 s -960 58428 480 58668 4 io_out[36]
port 135 nsew
rlabel metal3 s -960 19260 480 19500 4 io_out[37]
port 136 nsew
rlabel metal3 s 583520 139212 584960 139452 4 io_out[3]
port 137 nsew
rlabel metal3 s 583520 179060 584960 179300 4 io_out[4]
port 138 nsew
rlabel metal3 s 583520 218908 584960 219148 4 io_out[5]
port 139 nsew
rlabel metal3 s 583520 258756 584960 258996 4 io_out[6]
port 140 nsew
rlabel metal3 s 583520 311932 584960 312172 4 io_out[7]
port 141 nsew
rlabel metal3 s 583520 364972 584960 365212 4 io_out[8]
port 142 nsew
rlabel metal3 s 583520 418148 584960 418388 4 io_out[9]
port 143 nsew
rlabel metal2 s 125846 -960 125958 480 4 la_data_in[0]
port 144 nsew
rlabel metal2 s 480506 -960 480618 480 4 la_data_in[100]
port 145 nsew
rlabel metal2 s 484002 -960 484114 480 4 la_data_in[101]
port 146 nsew
rlabel metal2 s 487590 -960 487702 480 4 la_data_in[102]
port 147 nsew
rlabel metal2 s 491086 -960 491198 480 4 la_data_in[103]
port 148 nsew
rlabel metal2 s 494674 -960 494786 480 4 la_data_in[104]
port 149 nsew
rlabel metal2 s 498170 -960 498282 480 4 la_data_in[105]
port 150 nsew
rlabel metal2 s 501758 -960 501870 480 4 la_data_in[106]
port 151 nsew
rlabel metal2 s 505346 -960 505458 480 4 la_data_in[107]
port 152 nsew
rlabel metal2 s 508842 -960 508954 480 4 la_data_in[108]
port 153 nsew
rlabel metal2 s 512430 -960 512542 480 4 la_data_in[109]
port 154 nsew
rlabel metal2 s 161266 -960 161378 480 4 la_data_in[10]
port 155 nsew
rlabel metal2 s 515926 -960 516038 480 4 la_data_in[110]
port 156 nsew
rlabel metal2 s 519514 -960 519626 480 4 la_data_in[111]
port 157 nsew
rlabel metal2 s 523010 -960 523122 480 4 la_data_in[112]
port 158 nsew
rlabel metal2 s 526598 -960 526710 480 4 la_data_in[113]
port 159 nsew
rlabel metal2 s 530094 -960 530206 480 4 la_data_in[114]
port 160 nsew
rlabel metal2 s 533682 -960 533794 480 4 la_data_in[115]
port 161 nsew
rlabel metal2 s 537178 -960 537290 480 4 la_data_in[116]
port 162 nsew
rlabel metal2 s 540766 -960 540878 480 4 la_data_in[117]
port 163 nsew
rlabel metal2 s 544354 -960 544466 480 4 la_data_in[118]
port 164 nsew
rlabel metal2 s 547850 -960 547962 480 4 la_data_in[119]
port 165 nsew
rlabel metal2 s 164854 -960 164966 480 4 la_data_in[11]
port 166 nsew
rlabel metal2 s 551438 -960 551550 480 4 la_data_in[120]
port 167 nsew
rlabel metal2 s 554934 -960 555046 480 4 la_data_in[121]
port 168 nsew
rlabel metal2 s 558522 -960 558634 480 4 la_data_in[122]
port 169 nsew
rlabel metal2 s 562018 -960 562130 480 4 la_data_in[123]
port 170 nsew
rlabel metal2 s 565606 -960 565718 480 4 la_data_in[124]
port 171 nsew
rlabel metal2 s 569102 -960 569214 480 4 la_data_in[125]
port 172 nsew
rlabel metal2 s 572690 -960 572802 480 4 la_data_in[126]
port 173 nsew
rlabel metal2 s 576278 -960 576390 480 4 la_data_in[127]
port 174 nsew
rlabel metal2 s 168350 -960 168462 480 4 la_data_in[12]
port 175 nsew
rlabel metal2 s 171938 -960 172050 480 4 la_data_in[13]
port 176 nsew
rlabel metal2 s 175434 -960 175546 480 4 la_data_in[14]
port 177 nsew
rlabel metal2 s 179022 -960 179134 480 4 la_data_in[15]
port 178 nsew
rlabel metal2 s 182518 -960 182630 480 4 la_data_in[16]
port 179 nsew
rlabel metal2 s 186106 -960 186218 480 4 la_data_in[17]
port 180 nsew
rlabel metal2 s 189694 -960 189806 480 4 la_data_in[18]
port 181 nsew
rlabel metal2 s 193190 -960 193302 480 4 la_data_in[19]
port 182 nsew
rlabel metal2 s 129342 -960 129454 480 4 la_data_in[1]
port 183 nsew
rlabel metal2 s 196778 -960 196890 480 4 la_data_in[20]
port 184 nsew
rlabel metal2 s 200274 -960 200386 480 4 la_data_in[21]
port 185 nsew
rlabel metal2 s 203862 -960 203974 480 4 la_data_in[22]
port 186 nsew
rlabel metal2 s 207358 -960 207470 480 4 la_data_in[23]
port 187 nsew
rlabel metal2 s 210946 -960 211058 480 4 la_data_in[24]
port 188 nsew
rlabel metal2 s 214442 -960 214554 480 4 la_data_in[25]
port 189 nsew
rlabel metal2 s 218030 -960 218142 480 4 la_data_in[26]
port 190 nsew
rlabel metal2 s 221526 -960 221638 480 4 la_data_in[27]
port 191 nsew
rlabel metal2 s 225114 -960 225226 480 4 la_data_in[28]
port 192 nsew
rlabel metal2 s 228702 -960 228814 480 4 la_data_in[29]
port 193 nsew
rlabel metal2 s 132930 -960 133042 480 4 la_data_in[2]
port 194 nsew
rlabel metal2 s 232198 -960 232310 480 4 la_data_in[30]
port 195 nsew
rlabel metal2 s 235786 -960 235898 480 4 la_data_in[31]
port 196 nsew
rlabel metal2 s 239282 -960 239394 480 4 la_data_in[32]
port 197 nsew
rlabel metal2 s 242870 -960 242982 480 4 la_data_in[33]
port 198 nsew
rlabel metal2 s 246366 -960 246478 480 4 la_data_in[34]
port 199 nsew
rlabel metal2 s 249954 -960 250066 480 4 la_data_in[35]
port 200 nsew
rlabel metal2 s 253450 -960 253562 480 4 la_data_in[36]
port 201 nsew
rlabel metal2 s 257038 -960 257150 480 4 la_data_in[37]
port 202 nsew
rlabel metal2 s 260626 -960 260738 480 4 la_data_in[38]
port 203 nsew
rlabel metal2 s 264122 -960 264234 480 4 la_data_in[39]
port 204 nsew
rlabel metal2 s 136426 -960 136538 480 4 la_data_in[3]
port 205 nsew
rlabel metal2 s 267710 -960 267822 480 4 la_data_in[40]
port 206 nsew
rlabel metal2 s 271206 -960 271318 480 4 la_data_in[41]
port 207 nsew
rlabel metal2 s 274794 -960 274906 480 4 la_data_in[42]
port 208 nsew
rlabel metal2 s 278290 -960 278402 480 4 la_data_in[43]
port 209 nsew
rlabel metal2 s 281878 -960 281990 480 4 la_data_in[44]
port 210 nsew
rlabel metal2 s 285374 -960 285486 480 4 la_data_in[45]
port 211 nsew
rlabel metal2 s 288962 -960 289074 480 4 la_data_in[46]
port 212 nsew
rlabel metal2 s 292550 -960 292662 480 4 la_data_in[47]
port 213 nsew
rlabel metal2 s 296046 -960 296158 480 4 la_data_in[48]
port 214 nsew
rlabel metal2 s 299634 -960 299746 480 4 la_data_in[49]
port 215 nsew
rlabel metal2 s 140014 -960 140126 480 4 la_data_in[4]
port 216 nsew
rlabel metal2 s 303130 -960 303242 480 4 la_data_in[50]
port 217 nsew
rlabel metal2 s 306718 -960 306830 480 4 la_data_in[51]
port 218 nsew
rlabel metal2 s 310214 -960 310326 480 4 la_data_in[52]
port 219 nsew
rlabel metal2 s 313802 -960 313914 480 4 la_data_in[53]
port 220 nsew
rlabel metal2 s 317298 -960 317410 480 4 la_data_in[54]
port 221 nsew
rlabel metal2 s 320886 -960 320998 480 4 la_data_in[55]
port 222 nsew
rlabel metal2 s 324382 -960 324494 480 4 la_data_in[56]
port 223 nsew
rlabel metal2 s 327970 -960 328082 480 4 la_data_in[57]
port 224 nsew
rlabel metal2 s 331558 -960 331670 480 4 la_data_in[58]
port 225 nsew
rlabel metal2 s 335054 -960 335166 480 4 la_data_in[59]
port 226 nsew
rlabel metal2 s 143510 -960 143622 480 4 la_data_in[5]
port 227 nsew
rlabel metal2 s 338642 -960 338754 480 4 la_data_in[60]
port 228 nsew
rlabel metal2 s 342138 -960 342250 480 4 la_data_in[61]
port 229 nsew
rlabel metal2 s 345726 -960 345838 480 4 la_data_in[62]
port 230 nsew
rlabel metal2 s 349222 -960 349334 480 4 la_data_in[63]
port 231 nsew
rlabel metal2 s 352810 -960 352922 480 4 la_data_in[64]
port 232 nsew
rlabel metal2 s 356306 -960 356418 480 4 la_data_in[65]
port 233 nsew
rlabel metal2 s 359894 -960 360006 480 4 la_data_in[66]
port 234 nsew
rlabel metal2 s 363482 -960 363594 480 4 la_data_in[67]
port 235 nsew
rlabel metal2 s 366978 -960 367090 480 4 la_data_in[68]
port 236 nsew
rlabel metal2 s 370566 -960 370678 480 4 la_data_in[69]
port 237 nsew
rlabel metal2 s 147098 -960 147210 480 4 la_data_in[6]
port 238 nsew
rlabel metal2 s 374062 -960 374174 480 4 la_data_in[70]
port 239 nsew
rlabel metal2 s 377650 -960 377762 480 4 la_data_in[71]
port 240 nsew
rlabel metal2 s 381146 -960 381258 480 4 la_data_in[72]
port 241 nsew
rlabel metal2 s 384734 -960 384846 480 4 la_data_in[73]
port 242 nsew
rlabel metal2 s 388230 -960 388342 480 4 la_data_in[74]
port 243 nsew
rlabel metal2 s 391818 -960 391930 480 4 la_data_in[75]
port 244 nsew
rlabel metal2 s 395314 -960 395426 480 4 la_data_in[76]
port 245 nsew
rlabel metal2 s 398902 -960 399014 480 4 la_data_in[77]
port 246 nsew
rlabel metal2 s 402490 -960 402602 480 4 la_data_in[78]
port 247 nsew
rlabel metal2 s 405986 -960 406098 480 4 la_data_in[79]
port 248 nsew
rlabel metal2 s 150594 -960 150706 480 4 la_data_in[7]
port 249 nsew
rlabel metal2 s 409574 -960 409686 480 4 la_data_in[80]
port 250 nsew
rlabel metal2 s 413070 -960 413182 480 4 la_data_in[81]
port 251 nsew
rlabel metal2 s 416658 -960 416770 480 4 la_data_in[82]
port 252 nsew
rlabel metal2 s 420154 -960 420266 480 4 la_data_in[83]
port 253 nsew
rlabel metal2 s 423742 -960 423854 480 4 la_data_in[84]
port 254 nsew
rlabel metal2 s 427238 -960 427350 480 4 la_data_in[85]
port 255 nsew
rlabel metal2 s 430826 -960 430938 480 4 la_data_in[86]
port 256 nsew
rlabel metal2 s 434414 -960 434526 480 4 la_data_in[87]
port 257 nsew
rlabel metal2 s 437910 -960 438022 480 4 la_data_in[88]
port 258 nsew
rlabel metal2 s 441498 -960 441610 480 4 la_data_in[89]
port 259 nsew
rlabel metal2 s 154182 -960 154294 480 4 la_data_in[8]
port 260 nsew
rlabel metal2 s 444994 -960 445106 480 4 la_data_in[90]
port 261 nsew
rlabel metal2 s 448582 -960 448694 480 4 la_data_in[91]
port 262 nsew
rlabel metal2 s 452078 -960 452190 480 4 la_data_in[92]
port 263 nsew
rlabel metal2 s 455666 -960 455778 480 4 la_data_in[93]
port 264 nsew
rlabel metal2 s 459162 -960 459274 480 4 la_data_in[94]
port 265 nsew
rlabel metal2 s 462750 -960 462862 480 4 la_data_in[95]
port 266 nsew
rlabel metal2 s 466246 -960 466358 480 4 la_data_in[96]
port 267 nsew
rlabel metal2 s 469834 -960 469946 480 4 la_data_in[97]
port 268 nsew
rlabel metal2 s 473422 -960 473534 480 4 la_data_in[98]
port 269 nsew
rlabel metal2 s 476918 -960 477030 480 4 la_data_in[99]
port 270 nsew
rlabel metal2 s 157770 -960 157882 480 4 la_data_in[9]
port 271 nsew
rlabel metal2 s 126950 -960 127062 480 4 la_data_out[0]
port 272 nsew
rlabel metal2 s 481702 -960 481814 480 4 la_data_out[100]
port 273 nsew
rlabel metal2 s 485198 -960 485310 480 4 la_data_out[101]
port 274 nsew
rlabel metal2 s 488786 -960 488898 480 4 la_data_out[102]
port 275 nsew
rlabel metal2 s 492282 -960 492394 480 4 la_data_out[103]
port 276 nsew
rlabel metal2 s 495870 -960 495982 480 4 la_data_out[104]
port 277 nsew
rlabel metal2 s 499366 -960 499478 480 4 la_data_out[105]
port 278 nsew
rlabel metal2 s 502954 -960 503066 480 4 la_data_out[106]
port 279 nsew
rlabel metal2 s 506450 -960 506562 480 4 la_data_out[107]
port 280 nsew
rlabel metal2 s 510038 -960 510150 480 4 la_data_out[108]
port 281 nsew
rlabel metal2 s 513534 -960 513646 480 4 la_data_out[109]
port 282 nsew
rlabel metal2 s 162462 -960 162574 480 4 la_data_out[10]
port 283 nsew
rlabel metal2 s 517122 -960 517234 480 4 la_data_out[110]
port 284 nsew
rlabel metal2 s 520710 -960 520822 480 4 la_data_out[111]
port 285 nsew
rlabel metal2 s 524206 -960 524318 480 4 la_data_out[112]
port 286 nsew
rlabel metal2 s 527794 -960 527906 480 4 la_data_out[113]
port 287 nsew
rlabel metal2 s 531290 -960 531402 480 4 la_data_out[114]
port 288 nsew
rlabel metal2 s 534878 -960 534990 480 4 la_data_out[115]
port 289 nsew
rlabel metal2 s 538374 -960 538486 480 4 la_data_out[116]
port 290 nsew
rlabel metal2 s 541962 -960 542074 480 4 la_data_out[117]
port 291 nsew
rlabel metal2 s 545458 -960 545570 480 4 la_data_out[118]
port 292 nsew
rlabel metal2 s 549046 -960 549158 480 4 la_data_out[119]
port 293 nsew
rlabel metal2 s 166050 -960 166162 480 4 la_data_out[11]
port 294 nsew
rlabel metal2 s 552634 -960 552746 480 4 la_data_out[120]
port 295 nsew
rlabel metal2 s 556130 -960 556242 480 4 la_data_out[121]
port 296 nsew
rlabel metal2 s 559718 -960 559830 480 4 la_data_out[122]
port 297 nsew
rlabel metal2 s 563214 -960 563326 480 4 la_data_out[123]
port 298 nsew
rlabel metal2 s 566802 -960 566914 480 4 la_data_out[124]
port 299 nsew
rlabel metal2 s 570298 -960 570410 480 4 la_data_out[125]
port 300 nsew
rlabel metal2 s 573886 -960 573998 480 4 la_data_out[126]
port 301 nsew
rlabel metal2 s 577382 -960 577494 480 4 la_data_out[127]
port 302 nsew
rlabel metal2 s 169546 -960 169658 480 4 la_data_out[12]
port 303 nsew
rlabel metal2 s 173134 -960 173246 480 4 la_data_out[13]
port 304 nsew
rlabel metal2 s 176630 -960 176742 480 4 la_data_out[14]
port 305 nsew
rlabel metal2 s 180218 -960 180330 480 4 la_data_out[15]
port 306 nsew
rlabel metal2 s 183714 -960 183826 480 4 la_data_out[16]
port 307 nsew
rlabel metal2 s 187302 -960 187414 480 4 la_data_out[17]
port 308 nsew
rlabel metal2 s 190798 -960 190910 480 4 la_data_out[18]
port 309 nsew
rlabel metal2 s 194386 -960 194498 480 4 la_data_out[19]
port 310 nsew
rlabel metal2 s 130538 -960 130650 480 4 la_data_out[1]
port 311 nsew
rlabel metal2 s 197882 -960 197994 480 4 la_data_out[20]
port 312 nsew
rlabel metal2 s 201470 -960 201582 480 4 la_data_out[21]
port 313 nsew
rlabel metal2 s 205058 -960 205170 480 4 la_data_out[22]
port 314 nsew
rlabel metal2 s 208554 -960 208666 480 4 la_data_out[23]
port 315 nsew
rlabel metal2 s 212142 -960 212254 480 4 la_data_out[24]
port 316 nsew
rlabel metal2 s 215638 -960 215750 480 4 la_data_out[25]
port 317 nsew
rlabel metal2 s 219226 -960 219338 480 4 la_data_out[26]
port 318 nsew
rlabel metal2 s 222722 -960 222834 480 4 la_data_out[27]
port 319 nsew
rlabel metal2 s 226310 -960 226422 480 4 la_data_out[28]
port 320 nsew
rlabel metal2 s 229806 -960 229918 480 4 la_data_out[29]
port 321 nsew
rlabel metal2 s 134126 -960 134238 480 4 la_data_out[2]
port 322 nsew
rlabel metal2 s 233394 -960 233506 480 4 la_data_out[30]
port 323 nsew
rlabel metal2 s 236982 -960 237094 480 4 la_data_out[31]
port 324 nsew
rlabel metal2 s 240478 -960 240590 480 4 la_data_out[32]
port 325 nsew
rlabel metal2 s 244066 -960 244178 480 4 la_data_out[33]
port 326 nsew
rlabel metal2 s 247562 -960 247674 480 4 la_data_out[34]
port 327 nsew
rlabel metal2 s 251150 -960 251262 480 4 la_data_out[35]
port 328 nsew
rlabel metal2 s 254646 -960 254758 480 4 la_data_out[36]
port 329 nsew
rlabel metal2 s 258234 -960 258346 480 4 la_data_out[37]
port 330 nsew
rlabel metal2 s 261730 -960 261842 480 4 la_data_out[38]
port 331 nsew
rlabel metal2 s 265318 -960 265430 480 4 la_data_out[39]
port 332 nsew
rlabel metal2 s 137622 -960 137734 480 4 la_data_out[3]
port 333 nsew
rlabel metal2 s 268814 -960 268926 480 4 la_data_out[40]
port 334 nsew
rlabel metal2 s 272402 -960 272514 480 4 la_data_out[41]
port 335 nsew
rlabel metal2 s 275990 -960 276102 480 4 la_data_out[42]
port 336 nsew
rlabel metal2 s 279486 -960 279598 480 4 la_data_out[43]
port 337 nsew
rlabel metal2 s 283074 -960 283186 480 4 la_data_out[44]
port 338 nsew
rlabel metal2 s 286570 -960 286682 480 4 la_data_out[45]
port 339 nsew
rlabel metal2 s 290158 -960 290270 480 4 la_data_out[46]
port 340 nsew
rlabel metal2 s 293654 -960 293766 480 4 la_data_out[47]
port 341 nsew
rlabel metal2 s 297242 -960 297354 480 4 la_data_out[48]
port 342 nsew
rlabel metal2 s 300738 -960 300850 480 4 la_data_out[49]
port 343 nsew
rlabel metal2 s 141210 -960 141322 480 4 la_data_out[4]
port 344 nsew
rlabel metal2 s 304326 -960 304438 480 4 la_data_out[50]
port 345 nsew
rlabel metal2 s 307914 -960 308026 480 4 la_data_out[51]
port 346 nsew
rlabel metal2 s 311410 -960 311522 480 4 la_data_out[52]
port 347 nsew
rlabel metal2 s 314998 -960 315110 480 4 la_data_out[53]
port 348 nsew
rlabel metal2 s 318494 -960 318606 480 4 la_data_out[54]
port 349 nsew
rlabel metal2 s 322082 -960 322194 480 4 la_data_out[55]
port 350 nsew
rlabel metal2 s 325578 -960 325690 480 4 la_data_out[56]
port 351 nsew
rlabel metal2 s 329166 -960 329278 480 4 la_data_out[57]
port 352 nsew
rlabel metal2 s 332662 -960 332774 480 4 la_data_out[58]
port 353 nsew
rlabel metal2 s 336250 -960 336362 480 4 la_data_out[59]
port 354 nsew
rlabel metal2 s 144706 -960 144818 480 4 la_data_out[5]
port 355 nsew
rlabel metal2 s 339838 -960 339950 480 4 la_data_out[60]
port 356 nsew
rlabel metal2 s 343334 -960 343446 480 4 la_data_out[61]
port 357 nsew
rlabel metal2 s 346922 -960 347034 480 4 la_data_out[62]
port 358 nsew
rlabel metal2 s 350418 -960 350530 480 4 la_data_out[63]
port 359 nsew
rlabel metal2 s 354006 -960 354118 480 4 la_data_out[64]
port 360 nsew
rlabel metal2 s 357502 -960 357614 480 4 la_data_out[65]
port 361 nsew
rlabel metal2 s 361090 -960 361202 480 4 la_data_out[66]
port 362 nsew
rlabel metal2 s 364586 -960 364698 480 4 la_data_out[67]
port 363 nsew
rlabel metal2 s 368174 -960 368286 480 4 la_data_out[68]
port 364 nsew
rlabel metal2 s 371670 -960 371782 480 4 la_data_out[69]
port 365 nsew
rlabel metal2 s 148294 -960 148406 480 4 la_data_out[6]
port 366 nsew
rlabel metal2 s 375258 -960 375370 480 4 la_data_out[70]
port 367 nsew
rlabel metal2 s 378846 -960 378958 480 4 la_data_out[71]
port 368 nsew
rlabel metal2 s 382342 -960 382454 480 4 la_data_out[72]
port 369 nsew
rlabel metal2 s 385930 -960 386042 480 4 la_data_out[73]
port 370 nsew
rlabel metal2 s 389426 -960 389538 480 4 la_data_out[74]
port 371 nsew
rlabel metal2 s 393014 -960 393126 480 4 la_data_out[75]
port 372 nsew
rlabel metal2 s 396510 -960 396622 480 4 la_data_out[76]
port 373 nsew
rlabel metal2 s 400098 -960 400210 480 4 la_data_out[77]
port 374 nsew
rlabel metal2 s 403594 -960 403706 480 4 la_data_out[78]
port 375 nsew
rlabel metal2 s 407182 -960 407294 480 4 la_data_out[79]
port 376 nsew
rlabel metal2 s 151790 -960 151902 480 4 la_data_out[7]
port 377 nsew
rlabel metal2 s 410770 -960 410882 480 4 la_data_out[80]
port 378 nsew
rlabel metal2 s 414266 -960 414378 480 4 la_data_out[81]
port 379 nsew
rlabel metal2 s 417854 -960 417966 480 4 la_data_out[82]
port 380 nsew
rlabel metal2 s 421350 -960 421462 480 4 la_data_out[83]
port 381 nsew
rlabel metal2 s 424938 -960 425050 480 4 la_data_out[84]
port 382 nsew
rlabel metal2 s 428434 -960 428546 480 4 la_data_out[85]
port 383 nsew
rlabel metal2 s 432022 -960 432134 480 4 la_data_out[86]
port 384 nsew
rlabel metal2 s 435518 -960 435630 480 4 la_data_out[87]
port 385 nsew
rlabel metal2 s 439106 -960 439218 480 4 la_data_out[88]
port 386 nsew
rlabel metal2 s 442602 -960 442714 480 4 la_data_out[89]
port 387 nsew
rlabel metal2 s 155378 -960 155490 480 4 la_data_out[8]
port 388 nsew
rlabel metal2 s 446190 -960 446302 480 4 la_data_out[90]
port 389 nsew
rlabel metal2 s 449778 -960 449890 480 4 la_data_out[91]
port 390 nsew
rlabel metal2 s 453274 -960 453386 480 4 la_data_out[92]
port 391 nsew
rlabel metal2 s 456862 -960 456974 480 4 la_data_out[93]
port 392 nsew
rlabel metal2 s 460358 -960 460470 480 4 la_data_out[94]
port 393 nsew
rlabel metal2 s 463946 -960 464058 480 4 la_data_out[95]
port 394 nsew
rlabel metal2 s 467442 -960 467554 480 4 la_data_out[96]
port 395 nsew
rlabel metal2 s 471030 -960 471142 480 4 la_data_out[97]
port 396 nsew
rlabel metal2 s 474526 -960 474638 480 4 la_data_out[98]
port 397 nsew
rlabel metal2 s 478114 -960 478226 480 4 la_data_out[99]
port 398 nsew
rlabel metal2 s 158874 -960 158986 480 4 la_data_out[9]
port 399 nsew
rlabel metal2 s 128146 -960 128258 480 4 la_oenb[0]
port 400 nsew
rlabel metal2 s 482806 -960 482918 480 4 la_oenb[100]
port 401 nsew
rlabel metal2 s 486394 -960 486506 480 4 la_oenb[101]
port 402 nsew
rlabel metal2 s 489890 -960 490002 480 4 la_oenb[102]
port 403 nsew
rlabel metal2 s 493478 -960 493590 480 4 la_oenb[103]
port 404 nsew
rlabel metal2 s 497066 -960 497178 480 4 la_oenb[104]
port 405 nsew
rlabel metal2 s 500562 -960 500674 480 4 la_oenb[105]
port 406 nsew
rlabel metal2 s 504150 -960 504262 480 4 la_oenb[106]
port 407 nsew
rlabel metal2 s 507646 -960 507758 480 4 la_oenb[107]
port 408 nsew
rlabel metal2 s 511234 -960 511346 480 4 la_oenb[108]
port 409 nsew
rlabel metal2 s 514730 -960 514842 480 4 la_oenb[109]
port 410 nsew
rlabel metal2 s 163658 -960 163770 480 4 la_oenb[10]
port 411 nsew
rlabel metal2 s 518318 -960 518430 480 4 la_oenb[110]
port 412 nsew
rlabel metal2 s 521814 -960 521926 480 4 la_oenb[111]
port 413 nsew
rlabel metal2 s 525402 -960 525514 480 4 la_oenb[112]
port 414 nsew
rlabel metal2 s 528990 -960 529102 480 4 la_oenb[113]
port 415 nsew
rlabel metal2 s 532486 -960 532598 480 4 la_oenb[114]
port 416 nsew
rlabel metal2 s 536074 -960 536186 480 4 la_oenb[115]
port 417 nsew
rlabel metal2 s 539570 -960 539682 480 4 la_oenb[116]
port 418 nsew
rlabel metal2 s 543158 -960 543270 480 4 la_oenb[117]
port 419 nsew
rlabel metal2 s 546654 -960 546766 480 4 la_oenb[118]
port 420 nsew
rlabel metal2 s 550242 -960 550354 480 4 la_oenb[119]
port 421 nsew
rlabel metal2 s 167154 -960 167266 480 4 la_oenb[11]
port 422 nsew
rlabel metal2 s 553738 -960 553850 480 4 la_oenb[120]
port 423 nsew
rlabel metal2 s 557326 -960 557438 480 4 la_oenb[121]
port 424 nsew
rlabel metal2 s 560822 -960 560934 480 4 la_oenb[122]
port 425 nsew
rlabel metal2 s 564410 -960 564522 480 4 la_oenb[123]
port 426 nsew
rlabel metal2 s 567998 -960 568110 480 4 la_oenb[124]
port 427 nsew
rlabel metal2 s 571494 -960 571606 480 4 la_oenb[125]
port 428 nsew
rlabel metal2 s 575082 -960 575194 480 4 la_oenb[126]
port 429 nsew
rlabel metal2 s 578578 -960 578690 480 4 la_oenb[127]
port 430 nsew
rlabel metal2 s 170742 -960 170854 480 4 la_oenb[12]
port 431 nsew
rlabel metal2 s 174238 -960 174350 480 4 la_oenb[13]
port 432 nsew
rlabel metal2 s 177826 -960 177938 480 4 la_oenb[14]
port 433 nsew
rlabel metal2 s 181414 -960 181526 480 4 la_oenb[15]
port 434 nsew
rlabel metal2 s 184910 -960 185022 480 4 la_oenb[16]
port 435 nsew
rlabel metal2 s 188498 -960 188610 480 4 la_oenb[17]
port 436 nsew
rlabel metal2 s 191994 -960 192106 480 4 la_oenb[18]
port 437 nsew
rlabel metal2 s 195582 -960 195694 480 4 la_oenb[19]
port 438 nsew
rlabel metal2 s 131734 -960 131846 480 4 la_oenb[1]
port 439 nsew
rlabel metal2 s 199078 -960 199190 480 4 la_oenb[20]
port 440 nsew
rlabel metal2 s 202666 -960 202778 480 4 la_oenb[21]
port 441 nsew
rlabel metal2 s 206162 -960 206274 480 4 la_oenb[22]
port 442 nsew
rlabel metal2 s 209750 -960 209862 480 4 la_oenb[23]
port 443 nsew
rlabel metal2 s 213338 -960 213450 480 4 la_oenb[24]
port 444 nsew
rlabel metal2 s 216834 -960 216946 480 4 la_oenb[25]
port 445 nsew
rlabel metal2 s 220422 -960 220534 480 4 la_oenb[26]
port 446 nsew
rlabel metal2 s 223918 -960 224030 480 4 la_oenb[27]
port 447 nsew
rlabel metal2 s 227506 -960 227618 480 4 la_oenb[28]
port 448 nsew
rlabel metal2 s 231002 -960 231114 480 4 la_oenb[29]
port 449 nsew
rlabel metal2 s 135230 -960 135342 480 4 la_oenb[2]
port 450 nsew
rlabel metal2 s 234590 -960 234702 480 4 la_oenb[30]
port 451 nsew
rlabel metal2 s 238086 -960 238198 480 4 la_oenb[31]
port 452 nsew
rlabel metal2 s 241674 -960 241786 480 4 la_oenb[32]
port 453 nsew
rlabel metal2 s 245170 -960 245282 480 4 la_oenb[33]
port 454 nsew
rlabel metal2 s 248758 -960 248870 480 4 la_oenb[34]
port 455 nsew
rlabel metal2 s 252346 -960 252458 480 4 la_oenb[35]
port 456 nsew
rlabel metal2 s 255842 -960 255954 480 4 la_oenb[36]
port 457 nsew
rlabel metal2 s 259430 -960 259542 480 4 la_oenb[37]
port 458 nsew
rlabel metal2 s 262926 -960 263038 480 4 la_oenb[38]
port 459 nsew
rlabel metal2 s 266514 -960 266626 480 4 la_oenb[39]
port 460 nsew
rlabel metal2 s 138818 -960 138930 480 4 la_oenb[3]
port 461 nsew
rlabel metal2 s 270010 -960 270122 480 4 la_oenb[40]
port 462 nsew
rlabel metal2 s 273598 -960 273710 480 4 la_oenb[41]
port 463 nsew
rlabel metal2 s 277094 -960 277206 480 4 la_oenb[42]
port 464 nsew
rlabel metal2 s 280682 -960 280794 480 4 la_oenb[43]
port 465 nsew
rlabel metal2 s 284270 -960 284382 480 4 la_oenb[44]
port 466 nsew
rlabel metal2 s 287766 -960 287878 480 4 la_oenb[45]
port 467 nsew
rlabel metal2 s 291354 -960 291466 480 4 la_oenb[46]
port 468 nsew
rlabel metal2 s 294850 -960 294962 480 4 la_oenb[47]
port 469 nsew
rlabel metal2 s 298438 -960 298550 480 4 la_oenb[48]
port 470 nsew
rlabel metal2 s 301934 -960 302046 480 4 la_oenb[49]
port 471 nsew
rlabel metal2 s 142406 -960 142518 480 4 la_oenb[4]
port 472 nsew
rlabel metal2 s 305522 -960 305634 480 4 la_oenb[50]
port 473 nsew
rlabel metal2 s 309018 -960 309130 480 4 la_oenb[51]
port 474 nsew
rlabel metal2 s 312606 -960 312718 480 4 la_oenb[52]
port 475 nsew
rlabel metal2 s 316194 -960 316306 480 4 la_oenb[53]
port 476 nsew
rlabel metal2 s 319690 -960 319802 480 4 la_oenb[54]
port 477 nsew
rlabel metal2 s 323278 -960 323390 480 4 la_oenb[55]
port 478 nsew
rlabel metal2 s 326774 -960 326886 480 4 la_oenb[56]
port 479 nsew
rlabel metal2 s 330362 -960 330474 480 4 la_oenb[57]
port 480 nsew
rlabel metal2 s 333858 -960 333970 480 4 la_oenb[58]
port 481 nsew
rlabel metal2 s 337446 -960 337558 480 4 la_oenb[59]
port 482 nsew
rlabel metal2 s 145902 -960 146014 480 4 la_oenb[5]
port 483 nsew
rlabel metal2 s 340942 -960 341054 480 4 la_oenb[60]
port 484 nsew
rlabel metal2 s 344530 -960 344642 480 4 la_oenb[61]
port 485 nsew
rlabel metal2 s 348026 -960 348138 480 4 la_oenb[62]
port 486 nsew
rlabel metal2 s 351614 -960 351726 480 4 la_oenb[63]
port 487 nsew
rlabel metal2 s 355202 -960 355314 480 4 la_oenb[64]
port 488 nsew
rlabel metal2 s 358698 -960 358810 480 4 la_oenb[65]
port 489 nsew
rlabel metal2 s 362286 -960 362398 480 4 la_oenb[66]
port 490 nsew
rlabel metal2 s 365782 -960 365894 480 4 la_oenb[67]
port 491 nsew
rlabel metal2 s 369370 -960 369482 480 4 la_oenb[68]
port 492 nsew
rlabel metal2 s 372866 -960 372978 480 4 la_oenb[69]
port 493 nsew
rlabel metal2 s 149490 -960 149602 480 4 la_oenb[6]
port 494 nsew
rlabel metal2 s 376454 -960 376566 480 4 la_oenb[70]
port 495 nsew
rlabel metal2 s 379950 -960 380062 480 4 la_oenb[71]
port 496 nsew
rlabel metal2 s 383538 -960 383650 480 4 la_oenb[72]
port 497 nsew
rlabel metal2 s 387126 -960 387238 480 4 la_oenb[73]
port 498 nsew
rlabel metal2 s 390622 -960 390734 480 4 la_oenb[74]
port 499 nsew
rlabel metal2 s 394210 -960 394322 480 4 la_oenb[75]
port 500 nsew
rlabel metal2 s 397706 -960 397818 480 4 la_oenb[76]
port 501 nsew
rlabel metal2 s 401294 -960 401406 480 4 la_oenb[77]
port 502 nsew
rlabel metal2 s 404790 -960 404902 480 4 la_oenb[78]
port 503 nsew
rlabel metal2 s 408378 -960 408490 480 4 la_oenb[79]
port 504 nsew
rlabel metal2 s 152986 -960 153098 480 4 la_oenb[7]
port 505 nsew
rlabel metal2 s 411874 -960 411986 480 4 la_oenb[80]
port 506 nsew
rlabel metal2 s 415462 -960 415574 480 4 la_oenb[81]
port 507 nsew
rlabel metal2 s 418958 -960 419070 480 4 la_oenb[82]
port 508 nsew
rlabel metal2 s 422546 -960 422658 480 4 la_oenb[83]
port 509 nsew
rlabel metal2 s 426134 -960 426246 480 4 la_oenb[84]
port 510 nsew
rlabel metal2 s 429630 -960 429742 480 4 la_oenb[85]
port 511 nsew
rlabel metal2 s 433218 -960 433330 480 4 la_oenb[86]
port 512 nsew
rlabel metal2 s 436714 -960 436826 480 4 la_oenb[87]
port 513 nsew
rlabel metal2 s 440302 -960 440414 480 4 la_oenb[88]
port 514 nsew
rlabel metal2 s 443798 -960 443910 480 4 la_oenb[89]
port 515 nsew
rlabel metal2 s 156574 -960 156686 480 4 la_oenb[8]
port 516 nsew
rlabel metal2 s 447386 -960 447498 480 4 la_oenb[90]
port 517 nsew
rlabel metal2 s 450882 -960 450994 480 4 la_oenb[91]
port 518 nsew
rlabel metal2 s 454470 -960 454582 480 4 la_oenb[92]
port 519 nsew
rlabel metal2 s 458058 -960 458170 480 4 la_oenb[93]
port 520 nsew
rlabel metal2 s 461554 -960 461666 480 4 la_oenb[94]
port 521 nsew
rlabel metal2 s 465142 -960 465254 480 4 la_oenb[95]
port 522 nsew
rlabel metal2 s 468638 -960 468750 480 4 la_oenb[96]
port 523 nsew
rlabel metal2 s 472226 -960 472338 480 4 la_oenb[97]
port 524 nsew
rlabel metal2 s 475722 -960 475834 480 4 la_oenb[98]
port 525 nsew
rlabel metal2 s 479310 -960 479422 480 4 la_oenb[99]
port 526 nsew
rlabel metal2 s 160070 -960 160182 480 4 la_oenb[9]
port 527 nsew
rlabel metal2 s 579774 -960 579886 480 4 user_clock2
port 528 nsew
rlabel metal2 s 580970 -960 581082 480 4 user_irq[0]
port 529 nsew
rlabel metal2 s 582166 -960 582278 480 4 user_irq[1]
port 530 nsew
rlabel metal2 s 583362 -960 583474 480 4 user_irq[2]
port 531 nsew
rlabel metal5 s -2006 -934 585930 -314 4 vccd1
port 532 nsew
rlabel metal5 s -2966 2866 586890 3486 4 vccd1
port 532 nsew
rlabel metal5 s -2966 38866 586890 39486 4 vccd1
port 532 nsew
rlabel metal5 s -2966 74866 586890 75486 4 vccd1
port 532 nsew
rlabel metal5 s -2966 110866 586890 111486 4 vccd1
port 532 nsew
rlabel metal5 s -2966 146866 586890 147486 4 vccd1
port 532 nsew
rlabel metal5 s -2966 182866 586890 183486 4 vccd1
port 532 nsew
rlabel metal5 s -2966 218866 586890 219486 4 vccd1
port 532 nsew
rlabel metal5 s -2966 254866 586890 255486 4 vccd1
port 532 nsew
rlabel metal5 s -2966 290866 586890 291486 4 vccd1
port 532 nsew
rlabel metal5 s -2966 326866 586890 327486 4 vccd1
port 532 nsew
rlabel metal5 s -2966 362866 586890 363486 4 vccd1
port 532 nsew
rlabel metal5 s -2966 398866 586890 399486 4 vccd1
port 532 nsew
rlabel metal5 s -2966 434866 586890 435486 4 vccd1
port 532 nsew
rlabel metal5 s -2966 470866 586890 471486 4 vccd1
port 532 nsew
rlabel metal5 s -2966 506866 586890 507486 4 vccd1
port 532 nsew
rlabel metal5 s -2966 542866 586890 543486 4 vccd1
port 532 nsew
rlabel metal5 s -2966 578866 586890 579486 4 vccd1
port 532 nsew
rlabel metal5 s -2966 614866 586890 615486 4 vccd1
port 532 nsew
rlabel metal5 s -2966 650866 586890 651486 4 vccd1
port 532 nsew
rlabel metal5 s -2966 686866 586890 687486 4 vccd1
port 532 nsew
rlabel metal5 s -2006 704250 585930 704870 4 vccd1
port 532 nsew
rlabel metal4 s 253794 -1894 254414 336000 4 vccd1
port 532 nsew
rlabel metal4 s 289794 -1894 290414 336000 4 vccd1
port 532 nsew
rlabel metal4 s 325794 -1894 326414 336000 4 vccd1
port 532 nsew
rlabel metal4 s 361794 -1894 362414 336000 4 vccd1
port 532 nsew
rlabel metal4 s -2006 -934 -1386 704870 4 vccd1
port 532 nsew
rlabel metal4 s 585310 -934 585930 704870 4 vccd1
port 532 nsew
rlabel metal4 s 1794 -1894 2414 705830 4 vccd1
port 532 nsew
rlabel metal4 s 37794 -1894 38414 705830 4 vccd1
port 532 nsew
rlabel metal4 s 73794 -1894 74414 705830 4 vccd1
port 532 nsew
rlabel metal4 s 109794 -1894 110414 705830 4 vccd1
port 532 nsew
rlabel metal4 s 145794 -1894 146414 705830 4 vccd1
port 532 nsew
rlabel metal4 s 181794 -1894 182414 705830 4 vccd1
port 532 nsew
rlabel metal4 s 217794 -1894 218414 705830 4 vccd1
port 532 nsew
rlabel metal4 s 253794 489603 254414 705830 4 vccd1
port 532 nsew
rlabel metal4 s 289794 489603 290414 705830 4 vccd1
port 532 nsew
rlabel metal4 s 325794 489603 326414 705830 4 vccd1
port 532 nsew
rlabel metal4 s 361794 489603 362414 705830 4 vccd1
port 532 nsew
rlabel metal4 s 397794 -1894 398414 705830 4 vccd1
port 532 nsew
rlabel metal4 s 433794 -1894 434414 705830 4 vccd1
port 532 nsew
rlabel metal4 s 469794 -1894 470414 705830 4 vccd1
port 532 nsew
rlabel metal4 s 505794 -1894 506414 705830 4 vccd1
port 532 nsew
rlabel metal4 s 541794 -1894 542414 705830 4 vccd1
port 532 nsew
rlabel metal4 s 577794 -1894 578414 705830 4 vccd1
port 532 nsew
rlabel metal5 s -3926 -2854 587850 -2234 4 vccd2
port 533 nsew
rlabel metal5 s -4886 6586 588810 7206 4 vccd2
port 533 nsew
rlabel metal5 s -4886 42586 588810 43206 4 vccd2
port 533 nsew
rlabel metal5 s -4886 78586 588810 79206 4 vccd2
port 533 nsew
rlabel metal5 s -4886 114586 588810 115206 4 vccd2
port 533 nsew
rlabel metal5 s -4886 150586 588810 151206 4 vccd2
port 533 nsew
rlabel metal5 s -4886 186586 588810 187206 4 vccd2
port 533 nsew
rlabel metal5 s -4886 222586 588810 223206 4 vccd2
port 533 nsew
rlabel metal5 s -4886 258586 588810 259206 4 vccd2
port 533 nsew
rlabel metal5 s -4886 294586 588810 295206 4 vccd2
port 533 nsew
rlabel metal5 s -4886 330586 588810 331206 4 vccd2
port 533 nsew
rlabel metal5 s -4886 366586 588810 367206 4 vccd2
port 533 nsew
rlabel metal5 s -4886 402586 588810 403206 4 vccd2
port 533 nsew
rlabel metal5 s -4886 438586 588810 439206 4 vccd2
port 533 nsew
rlabel metal5 s -4886 474586 588810 475206 4 vccd2
port 533 nsew
rlabel metal5 s -4886 510586 588810 511206 4 vccd2
port 533 nsew
rlabel metal5 s -4886 546586 588810 547206 4 vccd2
port 533 nsew
rlabel metal5 s -4886 582586 588810 583206 4 vccd2
port 533 nsew
rlabel metal5 s -4886 618586 588810 619206 4 vccd2
port 533 nsew
rlabel metal5 s -4886 654586 588810 655206 4 vccd2
port 533 nsew
rlabel metal5 s -4886 690586 588810 691206 4 vccd2
port 533 nsew
rlabel metal5 s -3926 706170 587850 706790 4 vccd2
port 533 nsew
rlabel metal4 s 257514 -3814 258134 336000 4 vccd2
port 533 nsew
rlabel metal4 s 293514 -3814 294134 336000 4 vccd2
port 533 nsew
rlabel metal4 s 329514 -3814 330134 336000 4 vccd2
port 533 nsew
rlabel metal4 s 365514 -3814 366134 336000 4 vccd2
port 533 nsew
rlabel metal4 s -3926 -2854 -3306 706790 4 vccd2
port 533 nsew
rlabel metal4 s 587230 -2854 587850 706790 4 vccd2
port 533 nsew
rlabel metal4 s 5514 -3814 6134 707750 4 vccd2
port 533 nsew
rlabel metal4 s 41514 -3814 42134 707750 4 vccd2
port 533 nsew
rlabel metal4 s 77514 -3814 78134 707750 4 vccd2
port 533 nsew
rlabel metal4 s 113514 -3814 114134 707750 4 vccd2
port 533 nsew
rlabel metal4 s 149514 -3814 150134 707750 4 vccd2
port 533 nsew
rlabel metal4 s 185514 -3814 186134 707750 4 vccd2
port 533 nsew
rlabel metal4 s 221514 -3814 222134 707750 4 vccd2
port 533 nsew
rlabel metal4 s 257514 489603 258134 707750 4 vccd2
port 533 nsew
rlabel metal4 s 293514 489603 294134 707750 4 vccd2
port 533 nsew
rlabel metal4 s 329514 489603 330134 707750 4 vccd2
port 533 nsew
rlabel metal4 s 365514 489603 366134 707750 4 vccd2
port 533 nsew
rlabel metal4 s 401514 -3814 402134 707750 4 vccd2
port 533 nsew
rlabel metal4 s 437514 -3814 438134 707750 4 vccd2
port 533 nsew
rlabel metal4 s 473514 -3814 474134 707750 4 vccd2
port 533 nsew
rlabel metal4 s 509514 -3814 510134 707750 4 vccd2
port 533 nsew
rlabel metal4 s 545514 -3814 546134 707750 4 vccd2
port 533 nsew
rlabel metal4 s 581514 -3814 582134 707750 4 vccd2
port 533 nsew
rlabel metal5 s -5846 -4774 589770 -4154 4 vdda1
port 534 nsew
rlabel metal5 s -6806 10306 590730 10926 4 vdda1
port 534 nsew
rlabel metal5 s -6806 46306 590730 46926 4 vdda1
port 534 nsew
rlabel metal5 s -6806 82306 590730 82926 4 vdda1
port 534 nsew
rlabel metal5 s -6806 118306 590730 118926 4 vdda1
port 534 nsew
rlabel metal5 s -6806 154306 590730 154926 4 vdda1
port 534 nsew
rlabel metal5 s -6806 190306 590730 190926 4 vdda1
port 534 nsew
rlabel metal5 s -6806 226306 590730 226926 4 vdda1
port 534 nsew
rlabel metal5 s -6806 262306 590730 262926 4 vdda1
port 534 nsew
rlabel metal5 s -6806 298306 590730 298926 4 vdda1
port 534 nsew
rlabel metal5 s -6806 334306 590730 334926 4 vdda1
port 534 nsew
rlabel metal5 s -6806 370306 590730 370926 4 vdda1
port 534 nsew
rlabel metal5 s -6806 406306 590730 406926 4 vdda1
port 534 nsew
rlabel metal5 s -6806 442306 590730 442926 4 vdda1
port 534 nsew
rlabel metal5 s -6806 478306 590730 478926 4 vdda1
port 534 nsew
rlabel metal5 s -6806 514306 590730 514926 4 vdda1
port 534 nsew
rlabel metal5 s -6806 550306 590730 550926 4 vdda1
port 534 nsew
rlabel metal5 s -6806 586306 590730 586926 4 vdda1
port 534 nsew
rlabel metal5 s -6806 622306 590730 622926 4 vdda1
port 534 nsew
rlabel metal5 s -6806 658306 590730 658926 4 vdda1
port 534 nsew
rlabel metal5 s -6806 694306 590730 694926 4 vdda1
port 534 nsew
rlabel metal5 s -5846 708090 589770 708710 4 vdda1
port 534 nsew
rlabel metal4 s 261234 -5734 261854 336000 4 vdda1
port 534 nsew
rlabel metal4 s 297234 -5734 297854 336000 4 vdda1
port 534 nsew
rlabel metal4 s 333234 -5734 333854 336000 4 vdda1
port 534 nsew
rlabel metal4 s 369234 -5734 369854 336000 4 vdda1
port 534 nsew
rlabel metal4 s -5846 -4774 -5226 708710 4 vdda1
port 534 nsew
rlabel metal4 s 589150 -4774 589770 708710 4 vdda1
port 534 nsew
rlabel metal4 s 9234 -5734 9854 709670 4 vdda1
port 534 nsew
rlabel metal4 s 45234 -5734 45854 709670 4 vdda1
port 534 nsew
rlabel metal4 s 81234 -5734 81854 709670 4 vdda1
port 534 nsew
rlabel metal4 s 117234 -5734 117854 709670 4 vdda1
port 534 nsew
rlabel metal4 s 153234 -5734 153854 709670 4 vdda1
port 534 nsew
rlabel metal4 s 189234 -5734 189854 709670 4 vdda1
port 534 nsew
rlabel metal4 s 225234 -5734 225854 709670 4 vdda1
port 534 nsew
rlabel metal4 s 261234 489603 261854 709670 4 vdda1
port 534 nsew
rlabel metal4 s 297234 489603 297854 709670 4 vdda1
port 534 nsew
rlabel metal4 s 333234 489603 333854 709670 4 vdda1
port 534 nsew
rlabel metal4 s 369234 489603 369854 709670 4 vdda1
port 534 nsew
rlabel metal4 s 405234 -5734 405854 709670 4 vdda1
port 534 nsew
rlabel metal4 s 441234 -5734 441854 709670 4 vdda1
port 534 nsew
rlabel metal4 s 477234 -5734 477854 709670 4 vdda1
port 534 nsew
rlabel metal4 s 513234 -5734 513854 709670 4 vdda1
port 534 nsew
rlabel metal4 s 549234 -5734 549854 709670 4 vdda1
port 534 nsew
rlabel metal5 s -7766 -6694 591690 -6074 4 vdda2
port 535 nsew
rlabel metal5 s -8726 14026 592650 14646 4 vdda2
port 535 nsew
rlabel metal5 s -8726 50026 592650 50646 4 vdda2
port 535 nsew
rlabel metal5 s -8726 86026 592650 86646 4 vdda2
port 535 nsew
rlabel metal5 s -8726 122026 592650 122646 4 vdda2
port 535 nsew
rlabel metal5 s -8726 158026 592650 158646 4 vdda2
port 535 nsew
rlabel metal5 s -8726 194026 592650 194646 4 vdda2
port 535 nsew
rlabel metal5 s -8726 230026 592650 230646 4 vdda2
port 535 nsew
rlabel metal5 s -8726 266026 592650 266646 4 vdda2
port 535 nsew
rlabel metal5 s -8726 302026 592650 302646 4 vdda2
port 535 nsew
rlabel metal5 s -8726 338026 592650 338646 4 vdda2
port 535 nsew
rlabel metal5 s -8726 374026 592650 374646 4 vdda2
port 535 nsew
rlabel metal5 s -8726 410026 592650 410646 4 vdda2
port 535 nsew
rlabel metal5 s -8726 446026 592650 446646 4 vdda2
port 535 nsew
rlabel metal5 s -8726 482026 592650 482646 4 vdda2
port 535 nsew
rlabel metal5 s -8726 518026 592650 518646 4 vdda2
port 535 nsew
rlabel metal5 s -8726 554026 592650 554646 4 vdda2
port 535 nsew
rlabel metal5 s -8726 590026 592650 590646 4 vdda2
port 535 nsew
rlabel metal5 s -8726 626026 592650 626646 4 vdda2
port 535 nsew
rlabel metal5 s -8726 662026 592650 662646 4 vdda2
port 535 nsew
rlabel metal5 s -8726 698026 592650 698646 4 vdda2
port 535 nsew
rlabel metal5 s -7766 710010 591690 710630 4 vdda2
port 535 nsew
rlabel metal4 s 264954 -7654 265574 336000 4 vdda2
port 535 nsew
rlabel metal4 s 300954 -7654 301574 336000 4 vdda2
port 535 nsew
rlabel metal4 s 336954 -7654 337574 336000 4 vdda2
port 535 nsew
rlabel metal4 s 372954 -7654 373574 336000 4 vdda2
port 535 nsew
rlabel metal4 s -7766 -6694 -7146 710630 4 vdda2
port 535 nsew
rlabel metal4 s 591070 -6694 591690 710630 4 vdda2
port 535 nsew
rlabel metal4 s 12954 -7654 13574 711590 4 vdda2
port 535 nsew
rlabel metal4 s 48954 -7654 49574 711590 4 vdda2
port 535 nsew
rlabel metal4 s 84954 -7654 85574 711590 4 vdda2
port 535 nsew
rlabel metal4 s 120954 -7654 121574 711590 4 vdda2
port 535 nsew
rlabel metal4 s 156954 -7654 157574 711590 4 vdda2
port 535 nsew
rlabel metal4 s 192954 -7654 193574 711590 4 vdda2
port 535 nsew
rlabel metal4 s 228954 -7654 229574 711590 4 vdda2
port 535 nsew
rlabel metal4 s 264954 489603 265574 711590 4 vdda2
port 535 nsew
rlabel metal4 s 300954 489603 301574 711590 4 vdda2
port 535 nsew
rlabel metal4 s 336954 489603 337574 711590 4 vdda2
port 535 nsew
rlabel metal4 s 372954 489603 373574 711590 4 vdda2
port 535 nsew
rlabel metal4 s 408954 -7654 409574 711590 4 vdda2
port 535 nsew
rlabel metal4 s 444954 -7654 445574 711590 4 vdda2
port 535 nsew
rlabel metal4 s 480954 -7654 481574 711590 4 vdda2
port 535 nsew
rlabel metal4 s 516954 -7654 517574 711590 4 vdda2
port 535 nsew
rlabel metal4 s 552954 -7654 553574 711590 4 vdda2
port 535 nsew
rlabel metal5 s -6806 -5734 590730 -5114 4 vssa1
port 536 nsew
rlabel metal5 s -6806 28306 590730 28926 4 vssa1
port 536 nsew
rlabel metal5 s -6806 64306 590730 64926 4 vssa1
port 536 nsew
rlabel metal5 s -6806 100306 590730 100926 4 vssa1
port 536 nsew
rlabel metal5 s -6806 136306 590730 136926 4 vssa1
port 536 nsew
rlabel metal5 s -6806 172306 590730 172926 4 vssa1
port 536 nsew
rlabel metal5 s -6806 208306 590730 208926 4 vssa1
port 536 nsew
rlabel metal5 s -6806 244306 590730 244926 4 vssa1
port 536 nsew
rlabel metal5 s -6806 280306 590730 280926 4 vssa1
port 536 nsew
rlabel metal5 s -6806 316306 590730 316926 4 vssa1
port 536 nsew
rlabel metal5 s -6806 352306 590730 352926 4 vssa1
port 536 nsew
rlabel metal5 s -6806 388306 590730 388926 4 vssa1
port 536 nsew
rlabel metal5 s -6806 424306 590730 424926 4 vssa1
port 536 nsew
rlabel metal5 s -6806 460306 590730 460926 4 vssa1
port 536 nsew
rlabel metal5 s -6806 496306 590730 496926 4 vssa1
port 536 nsew
rlabel metal5 s -6806 532306 590730 532926 4 vssa1
port 536 nsew
rlabel metal5 s -6806 568306 590730 568926 4 vssa1
port 536 nsew
rlabel metal5 s -6806 604306 590730 604926 4 vssa1
port 536 nsew
rlabel metal5 s -6806 640306 590730 640926 4 vssa1
port 536 nsew
rlabel metal5 s -6806 676306 590730 676926 4 vssa1
port 536 nsew
rlabel metal5 s -6806 709050 590730 709670 4 vssa1
port 536 nsew
rlabel metal4 s 243234 -5734 243854 336000 4 vssa1
port 536 nsew
rlabel metal4 s 279234 -5734 279854 336000 4 vssa1
port 536 nsew
rlabel metal4 s 315234 -5734 315854 336000 4 vssa1
port 536 nsew
rlabel metal4 s 351234 -5734 351854 336000 4 vssa1
port 536 nsew
rlabel metal4 s -6806 -5734 -6186 709670 4 vssa1
port 536 nsew
rlabel metal4 s 27234 -5734 27854 709670 4 vssa1
port 536 nsew
rlabel metal4 s 63234 -5734 63854 709670 4 vssa1
port 536 nsew
rlabel metal4 s 99234 -5734 99854 709670 4 vssa1
port 536 nsew
rlabel metal4 s 135234 -5734 135854 709670 4 vssa1
port 536 nsew
rlabel metal4 s 171234 -5734 171854 709670 4 vssa1
port 536 nsew
rlabel metal4 s 207234 -5734 207854 709670 4 vssa1
port 536 nsew
rlabel metal4 s 243234 489603 243854 709670 4 vssa1
port 536 nsew
rlabel metal4 s 279234 489603 279854 709670 4 vssa1
port 536 nsew
rlabel metal4 s 315234 489603 315854 709670 4 vssa1
port 536 nsew
rlabel metal4 s 351234 489603 351854 709670 4 vssa1
port 536 nsew
rlabel metal4 s 387234 -5734 387854 709670 4 vssa1
port 536 nsew
rlabel metal4 s 423234 -5734 423854 709670 4 vssa1
port 536 nsew
rlabel metal4 s 459234 -5734 459854 709670 4 vssa1
port 536 nsew
rlabel metal4 s 495234 -5734 495854 709670 4 vssa1
port 536 nsew
rlabel metal4 s 531234 -5734 531854 709670 4 vssa1
port 536 nsew
rlabel metal4 s 567234 -5734 567854 709670 4 vssa1
port 536 nsew
rlabel metal4 s 590110 -5734 590730 709670 4 vssa1
port 536 nsew
rlabel metal5 s -8726 -7654 592650 -7034 4 vssa2
port 537 nsew
rlabel metal5 s -8726 32026 592650 32646 4 vssa2
port 537 nsew
rlabel metal5 s -8726 68026 592650 68646 4 vssa2
port 537 nsew
rlabel metal5 s -8726 104026 592650 104646 4 vssa2
port 537 nsew
rlabel metal5 s -8726 140026 592650 140646 4 vssa2
port 537 nsew
rlabel metal5 s -8726 176026 592650 176646 4 vssa2
port 537 nsew
rlabel metal5 s -8726 212026 592650 212646 4 vssa2
port 537 nsew
rlabel metal5 s -8726 248026 592650 248646 4 vssa2
port 537 nsew
rlabel metal5 s -8726 284026 592650 284646 4 vssa2
port 537 nsew
rlabel metal5 s -8726 320026 592650 320646 4 vssa2
port 537 nsew
rlabel metal5 s -8726 356026 592650 356646 4 vssa2
port 537 nsew
rlabel metal5 s -8726 392026 592650 392646 4 vssa2
port 537 nsew
rlabel metal5 s -8726 428026 592650 428646 4 vssa2
port 537 nsew
rlabel metal5 s -8726 464026 592650 464646 4 vssa2
port 537 nsew
rlabel metal5 s -8726 500026 592650 500646 4 vssa2
port 537 nsew
rlabel metal5 s -8726 536026 592650 536646 4 vssa2
port 537 nsew
rlabel metal5 s -8726 572026 592650 572646 4 vssa2
port 537 nsew
rlabel metal5 s -8726 608026 592650 608646 4 vssa2
port 537 nsew
rlabel metal5 s -8726 644026 592650 644646 4 vssa2
port 537 nsew
rlabel metal5 s -8726 680026 592650 680646 4 vssa2
port 537 nsew
rlabel metal5 s -8726 710970 592650 711590 4 vssa2
port 537 nsew
rlabel metal4 s 246954 -7654 247574 336000 4 vssa2
port 537 nsew
rlabel metal4 s 282954 -7654 283574 336000 4 vssa2
port 537 nsew
rlabel metal4 s 318954 -7654 319574 336000 4 vssa2
port 537 nsew
rlabel metal4 s 354954 -7654 355574 336000 4 vssa2
port 537 nsew
rlabel metal4 s -8726 -7654 -8106 711590 4 vssa2
port 537 nsew
rlabel metal4 s 30954 -7654 31574 711590 4 vssa2
port 537 nsew
rlabel metal4 s 66954 -7654 67574 711590 4 vssa2
port 537 nsew
rlabel metal4 s 102954 -7654 103574 711590 4 vssa2
port 537 nsew
rlabel metal4 s 138954 -7654 139574 711590 4 vssa2
port 537 nsew
rlabel metal4 s 174954 -7654 175574 711590 4 vssa2
port 537 nsew
rlabel metal4 s 210954 -7654 211574 711590 4 vssa2
port 537 nsew
rlabel metal4 s 246954 489603 247574 711590 4 vssa2
port 537 nsew
rlabel metal4 s 282954 489603 283574 711590 4 vssa2
port 537 nsew
rlabel metal4 s 318954 489603 319574 711590 4 vssa2
port 537 nsew
rlabel metal4 s 354954 489603 355574 711590 4 vssa2
port 537 nsew
rlabel metal4 s 390954 -7654 391574 711590 4 vssa2
port 537 nsew
rlabel metal4 s 426954 -7654 427574 711590 4 vssa2
port 537 nsew
rlabel metal4 s 462954 -7654 463574 711590 4 vssa2
port 537 nsew
rlabel metal4 s 498954 -7654 499574 711590 4 vssa2
port 537 nsew
rlabel metal4 s 534954 -7654 535574 711590 4 vssa2
port 537 nsew
rlabel metal4 s 570954 -7654 571574 711590 4 vssa2
port 537 nsew
rlabel metal4 s 592030 -7654 592650 711590 4 vssa2
port 537 nsew
rlabel metal5 s -2966 -1894 586890 -1274 4 vssd1
port 538 nsew
rlabel metal5 s -2966 20866 586890 21486 4 vssd1
port 538 nsew
rlabel metal5 s -2966 56866 586890 57486 4 vssd1
port 538 nsew
rlabel metal5 s -2966 92866 586890 93486 4 vssd1
port 538 nsew
rlabel metal5 s -2966 128866 586890 129486 4 vssd1
port 538 nsew
rlabel metal5 s -2966 164866 586890 165486 4 vssd1
port 538 nsew
rlabel metal5 s -2966 200866 586890 201486 4 vssd1
port 538 nsew
rlabel metal5 s -2966 236866 586890 237486 4 vssd1
port 538 nsew
rlabel metal5 s -2966 272866 586890 273486 4 vssd1
port 538 nsew
rlabel metal5 s -2966 308866 586890 309486 4 vssd1
port 538 nsew
rlabel metal5 s -2966 344866 586890 345486 4 vssd1
port 538 nsew
rlabel metal5 s -2966 380866 586890 381486 4 vssd1
port 538 nsew
rlabel metal5 s -2966 416866 586890 417486 4 vssd1
port 538 nsew
rlabel metal5 s -2966 452866 586890 453486 4 vssd1
port 538 nsew
rlabel metal5 s -2966 488866 586890 489486 4 vssd1
port 538 nsew
rlabel metal5 s -2966 524866 586890 525486 4 vssd1
port 538 nsew
rlabel metal5 s -2966 560866 586890 561486 4 vssd1
port 538 nsew
rlabel metal5 s -2966 596866 586890 597486 4 vssd1
port 538 nsew
rlabel metal5 s -2966 632866 586890 633486 4 vssd1
port 538 nsew
rlabel metal5 s -2966 668866 586890 669486 4 vssd1
port 538 nsew
rlabel metal5 s -2966 705210 586890 705830 4 vssd1
port 538 nsew
rlabel metal4 s 235794 -1894 236414 336000 4 vssd1
port 538 nsew
rlabel metal4 s 271794 -1894 272414 336000 4 vssd1
port 538 nsew
rlabel metal4 s 307794 -1894 308414 336000 4 vssd1
port 538 nsew
rlabel metal4 s 343794 -1894 344414 336000 4 vssd1
port 538 nsew
rlabel metal4 s 379794 -1894 380414 336000 4 vssd1
port 538 nsew
rlabel metal4 s -2966 -1894 -2346 705830 4 vssd1
port 538 nsew
rlabel metal4 s 19794 -1894 20414 705830 4 vssd1
port 538 nsew
rlabel metal4 s 55794 -1894 56414 705830 4 vssd1
port 538 nsew
rlabel metal4 s 91794 -1894 92414 705830 4 vssd1
port 538 nsew
rlabel metal4 s 127794 -1894 128414 705830 4 vssd1
port 538 nsew
rlabel metal4 s 163794 -1894 164414 705830 4 vssd1
port 538 nsew
rlabel metal4 s 199794 -1894 200414 705830 4 vssd1
port 538 nsew
rlabel metal4 s 235794 489603 236414 705830 4 vssd1
port 538 nsew
rlabel metal4 s 271794 489603 272414 705830 4 vssd1
port 538 nsew
rlabel metal4 s 307794 489603 308414 705830 4 vssd1
port 538 nsew
rlabel metal4 s 343794 489603 344414 705830 4 vssd1
port 538 nsew
rlabel metal4 s 379794 489603 380414 705830 4 vssd1
port 538 nsew
rlabel metal4 s 415794 -1894 416414 705830 4 vssd1
port 538 nsew
rlabel metal4 s 451794 -1894 452414 705830 4 vssd1
port 538 nsew
rlabel metal4 s 487794 -1894 488414 705830 4 vssd1
port 538 nsew
rlabel metal4 s 523794 -1894 524414 705830 4 vssd1
port 538 nsew
rlabel metal4 s 559794 -1894 560414 705830 4 vssd1
port 538 nsew
rlabel metal4 s 586270 -1894 586890 705830 4 vssd1
port 538 nsew
rlabel metal5 s -4886 -3814 588810 -3194 4 vssd2
port 539 nsew
rlabel metal5 s -4886 24586 588810 25206 4 vssd2
port 539 nsew
rlabel metal5 s -4886 60586 588810 61206 4 vssd2
port 539 nsew
rlabel metal5 s -4886 96586 588810 97206 4 vssd2
port 539 nsew
rlabel metal5 s -4886 132586 588810 133206 4 vssd2
port 539 nsew
rlabel metal5 s -4886 168586 588810 169206 4 vssd2
port 539 nsew
rlabel metal5 s -4886 204586 588810 205206 4 vssd2
port 539 nsew
rlabel metal5 s -4886 240586 588810 241206 4 vssd2
port 539 nsew
rlabel metal5 s -4886 276586 588810 277206 4 vssd2
port 539 nsew
rlabel metal5 s -4886 312586 588810 313206 4 vssd2
port 539 nsew
rlabel metal5 s -4886 348586 588810 349206 4 vssd2
port 539 nsew
rlabel metal5 s -4886 384586 588810 385206 4 vssd2
port 539 nsew
rlabel metal5 s -4886 420586 588810 421206 4 vssd2
port 539 nsew
rlabel metal5 s -4886 456586 588810 457206 4 vssd2
port 539 nsew
rlabel metal5 s -4886 492586 588810 493206 4 vssd2
port 539 nsew
rlabel metal5 s -4886 528586 588810 529206 4 vssd2
port 539 nsew
rlabel metal5 s -4886 564586 588810 565206 4 vssd2
port 539 nsew
rlabel metal5 s -4886 600586 588810 601206 4 vssd2
port 539 nsew
rlabel metal5 s -4886 636586 588810 637206 4 vssd2
port 539 nsew
rlabel metal5 s -4886 672586 588810 673206 4 vssd2
port 539 nsew
rlabel metal5 s -4886 707130 588810 707750 4 vssd2
port 539 nsew
rlabel metal4 s 239514 -3814 240134 336000 4 vssd2
port 539 nsew
rlabel metal4 s 275514 -3814 276134 336000 4 vssd2
port 539 nsew
rlabel metal4 s 311514 -3814 312134 336000 4 vssd2
port 539 nsew
rlabel metal4 s 347514 -3814 348134 336000 4 vssd2
port 539 nsew
rlabel metal4 s 383514 -3814 384134 336000 4 vssd2
port 539 nsew
rlabel metal4 s -4886 -3814 -4266 707750 4 vssd2
port 539 nsew
rlabel metal4 s 23514 -3814 24134 707750 4 vssd2
port 539 nsew
rlabel metal4 s 59514 -3814 60134 707750 4 vssd2
port 539 nsew
rlabel metal4 s 95514 -3814 96134 707750 4 vssd2
port 539 nsew
rlabel metal4 s 131514 -3814 132134 707750 4 vssd2
port 539 nsew
rlabel metal4 s 167514 -3814 168134 707750 4 vssd2
port 539 nsew
rlabel metal4 s 203514 -3814 204134 707750 4 vssd2
port 539 nsew
rlabel metal4 s 239514 489603 240134 707750 4 vssd2
port 539 nsew
rlabel metal4 s 275514 489603 276134 707750 4 vssd2
port 539 nsew
rlabel metal4 s 311514 489603 312134 707750 4 vssd2
port 539 nsew
rlabel metal4 s 347514 489603 348134 707750 4 vssd2
port 539 nsew
rlabel metal4 s 383514 489603 384134 707750 4 vssd2
port 539 nsew
rlabel metal4 s 419514 -3814 420134 707750 4 vssd2
port 539 nsew
rlabel metal4 s 455514 -3814 456134 707750 4 vssd2
port 539 nsew
rlabel metal4 s 491514 -3814 492134 707750 4 vssd2
port 539 nsew
rlabel metal4 s 527514 -3814 528134 707750 4 vssd2
port 539 nsew
rlabel metal4 s 563514 -3814 564134 707750 4 vssd2
port 539 nsew
rlabel metal4 s 588190 -3814 588810 707750 4 vssd2
port 539 nsew
rlabel metal2 s 542 -960 654 480 4 wb_clk_i
port 540 nsew
rlabel metal2 s 1646 -960 1758 480 4 wb_rst_i
port 541 nsew
rlabel metal2 s 2842 -960 2954 480 4 wbs_ack_o
port 542 nsew
rlabel metal2 s 7626 -960 7738 480 4 wbs_adr_i[0]
port 543 nsew
rlabel metal2 s 47830 -960 47942 480 4 wbs_adr_i[10]
port 544 nsew
rlabel metal2 s 51326 -960 51438 480 4 wbs_adr_i[11]
port 545 nsew
rlabel metal2 s 54914 -960 55026 480 4 wbs_adr_i[12]
port 546 nsew
rlabel metal2 s 58410 -960 58522 480 4 wbs_adr_i[13]
port 547 nsew
rlabel metal2 s 61998 -960 62110 480 4 wbs_adr_i[14]
port 548 nsew
rlabel metal2 s 65494 -960 65606 480 4 wbs_adr_i[15]
port 549 nsew
rlabel metal2 s 69082 -960 69194 480 4 wbs_adr_i[16]
port 550 nsew
rlabel metal2 s 72578 -960 72690 480 4 wbs_adr_i[17]
port 551 nsew
rlabel metal2 s 76166 -960 76278 480 4 wbs_adr_i[18]
port 552 nsew
rlabel metal2 s 79662 -960 79774 480 4 wbs_adr_i[19]
port 553 nsew
rlabel metal2 s 12318 -960 12430 480 4 wbs_adr_i[1]
port 554 nsew
rlabel metal2 s 83250 -960 83362 480 4 wbs_adr_i[20]
port 555 nsew
rlabel metal2 s 86838 -960 86950 480 4 wbs_adr_i[21]
port 556 nsew
rlabel metal2 s 90334 -960 90446 480 4 wbs_adr_i[22]
port 557 nsew
rlabel metal2 s 93922 -960 94034 480 4 wbs_adr_i[23]
port 558 nsew
rlabel metal2 s 97418 -960 97530 480 4 wbs_adr_i[24]
port 559 nsew
rlabel metal2 s 101006 -960 101118 480 4 wbs_adr_i[25]
port 560 nsew
rlabel metal2 s 104502 -960 104614 480 4 wbs_adr_i[26]
port 561 nsew
rlabel metal2 s 108090 -960 108202 480 4 wbs_adr_i[27]
port 562 nsew
rlabel metal2 s 111586 -960 111698 480 4 wbs_adr_i[28]
port 563 nsew
rlabel metal2 s 115174 -960 115286 480 4 wbs_adr_i[29]
port 564 nsew
rlabel metal2 s 17010 -960 17122 480 4 wbs_adr_i[2]
port 565 nsew
rlabel metal2 s 118762 -960 118874 480 4 wbs_adr_i[30]
port 566 nsew
rlabel metal2 s 122258 -960 122370 480 4 wbs_adr_i[31]
port 567 nsew
rlabel metal2 s 21794 -960 21906 480 4 wbs_adr_i[3]
port 568 nsew
rlabel metal2 s 26486 -960 26598 480 4 wbs_adr_i[4]
port 569 nsew
rlabel metal2 s 30074 -960 30186 480 4 wbs_adr_i[5]
port 570 nsew
rlabel metal2 s 33570 -960 33682 480 4 wbs_adr_i[6]
port 571 nsew
rlabel metal2 s 37158 -960 37270 480 4 wbs_adr_i[7]
port 572 nsew
rlabel metal2 s 40654 -960 40766 480 4 wbs_adr_i[8]
port 573 nsew
rlabel metal2 s 44242 -960 44354 480 4 wbs_adr_i[9]
port 574 nsew
rlabel metal2 s 4038 -960 4150 480 4 wbs_cyc_i
port 575 nsew
rlabel metal2 s 8730 -960 8842 480 4 wbs_dat_i[0]
port 576 nsew
rlabel metal2 s 48934 -960 49046 480 4 wbs_dat_i[10]
port 577 nsew
rlabel metal2 s 52522 -960 52634 480 4 wbs_dat_i[11]
port 578 nsew
rlabel metal2 s 56018 -960 56130 480 4 wbs_dat_i[12]
port 579 nsew
rlabel metal2 s 59606 -960 59718 480 4 wbs_dat_i[13]
port 580 nsew
rlabel metal2 s 63194 -960 63306 480 4 wbs_dat_i[14]
port 581 nsew
rlabel metal2 s 66690 -960 66802 480 4 wbs_dat_i[15]
port 582 nsew
rlabel metal2 s 70278 -960 70390 480 4 wbs_dat_i[16]
port 583 nsew
rlabel metal2 s 73774 -960 73886 480 4 wbs_dat_i[17]
port 584 nsew
rlabel metal2 s 77362 -960 77474 480 4 wbs_dat_i[18]
port 585 nsew
rlabel metal2 s 80858 -960 80970 480 4 wbs_dat_i[19]
port 586 nsew
rlabel metal2 s 13514 -960 13626 480 4 wbs_dat_i[1]
port 587 nsew
rlabel metal2 s 84446 -960 84558 480 4 wbs_dat_i[20]
port 588 nsew
rlabel metal2 s 87942 -960 88054 480 4 wbs_dat_i[21]
port 589 nsew
rlabel metal2 s 91530 -960 91642 480 4 wbs_dat_i[22]
port 590 nsew
rlabel metal2 s 95118 -960 95230 480 4 wbs_dat_i[23]
port 591 nsew
rlabel metal2 s 98614 -960 98726 480 4 wbs_dat_i[24]
port 592 nsew
rlabel metal2 s 102202 -960 102314 480 4 wbs_dat_i[25]
port 593 nsew
rlabel metal2 s 105698 -960 105810 480 4 wbs_dat_i[26]
port 594 nsew
rlabel metal2 s 109286 -960 109398 480 4 wbs_dat_i[27]
port 595 nsew
rlabel metal2 s 112782 -960 112894 480 4 wbs_dat_i[28]
port 596 nsew
rlabel metal2 s 116370 -960 116482 480 4 wbs_dat_i[29]
port 597 nsew
rlabel metal2 s 18206 -960 18318 480 4 wbs_dat_i[2]
port 598 nsew
rlabel metal2 s 119866 -960 119978 480 4 wbs_dat_i[30]
port 599 nsew
rlabel metal2 s 123454 -960 123566 480 4 wbs_dat_i[31]
port 600 nsew
rlabel metal2 s 22990 -960 23102 480 4 wbs_dat_i[3]
port 601 nsew
rlabel metal2 s 27682 -960 27794 480 4 wbs_dat_i[4]
port 602 nsew
rlabel metal2 s 31270 -960 31382 480 4 wbs_dat_i[5]
port 603 nsew
rlabel metal2 s 34766 -960 34878 480 4 wbs_dat_i[6]
port 604 nsew
rlabel metal2 s 38354 -960 38466 480 4 wbs_dat_i[7]
port 605 nsew
rlabel metal2 s 41850 -960 41962 480 4 wbs_dat_i[8]
port 606 nsew
rlabel metal2 s 45438 -960 45550 480 4 wbs_dat_i[9]
port 607 nsew
rlabel metal2 s 9926 -960 10038 480 4 wbs_dat_o[0]
port 608 nsew
rlabel metal2 s 50130 -960 50242 480 4 wbs_dat_o[10]
port 609 nsew
rlabel metal2 s 53718 -960 53830 480 4 wbs_dat_o[11]
port 610 nsew
rlabel metal2 s 57214 -960 57326 480 4 wbs_dat_o[12]
port 611 nsew
rlabel metal2 s 60802 -960 60914 480 4 wbs_dat_o[13]
port 612 nsew
rlabel metal2 s 64298 -960 64410 480 4 wbs_dat_o[14]
port 613 nsew
rlabel metal2 s 67886 -960 67998 480 4 wbs_dat_o[15]
port 614 nsew
rlabel metal2 s 71474 -960 71586 480 4 wbs_dat_o[16]
port 615 nsew
rlabel metal2 s 74970 -960 75082 480 4 wbs_dat_o[17]
port 616 nsew
rlabel metal2 s 78558 -960 78670 480 4 wbs_dat_o[18]
port 617 nsew
rlabel metal2 s 82054 -960 82166 480 4 wbs_dat_o[19]
port 618 nsew
rlabel metal2 s 14710 -960 14822 480 4 wbs_dat_o[1]
port 619 nsew
rlabel metal2 s 85642 -960 85754 480 4 wbs_dat_o[20]
port 620 nsew
rlabel metal2 s 89138 -960 89250 480 4 wbs_dat_o[21]
port 621 nsew
rlabel metal2 s 92726 -960 92838 480 4 wbs_dat_o[22]
port 622 nsew
rlabel metal2 s 96222 -960 96334 480 4 wbs_dat_o[23]
port 623 nsew
rlabel metal2 s 99810 -960 99922 480 4 wbs_dat_o[24]
port 624 nsew
rlabel metal2 s 103306 -960 103418 480 4 wbs_dat_o[25]
port 625 nsew
rlabel metal2 s 106894 -960 107006 480 4 wbs_dat_o[26]
port 626 nsew
rlabel metal2 s 110482 -960 110594 480 4 wbs_dat_o[27]
port 627 nsew
rlabel metal2 s 113978 -960 114090 480 4 wbs_dat_o[28]
port 628 nsew
rlabel metal2 s 117566 -960 117678 480 4 wbs_dat_o[29]
port 629 nsew
rlabel metal2 s 19402 -960 19514 480 4 wbs_dat_o[2]
port 630 nsew
rlabel metal2 s 121062 -960 121174 480 4 wbs_dat_o[30]
port 631 nsew
rlabel metal2 s 124650 -960 124762 480 4 wbs_dat_o[31]
port 632 nsew
rlabel metal2 s 24186 -960 24298 480 4 wbs_dat_o[3]
port 633 nsew
rlabel metal2 s 28878 -960 28990 480 4 wbs_dat_o[4]
port 634 nsew
rlabel metal2 s 32374 -960 32486 480 4 wbs_dat_o[5]
port 635 nsew
rlabel metal2 s 35962 -960 36074 480 4 wbs_dat_o[6]
port 636 nsew
rlabel metal2 s 39550 -960 39662 480 4 wbs_dat_o[7]
port 637 nsew
rlabel metal2 s 43046 -960 43158 480 4 wbs_dat_o[8]
port 638 nsew
rlabel metal2 s 46634 -960 46746 480 4 wbs_dat_o[9]
port 639 nsew
rlabel metal2 s 11122 -960 11234 480 4 wbs_sel_i[0]
port 640 nsew
rlabel metal2 s 15906 -960 16018 480 4 wbs_sel_i[1]
port 641 nsew
rlabel metal2 s 20598 -960 20710 480 4 wbs_sel_i[2]
port 642 nsew
rlabel metal2 s 25290 -960 25402 480 4 wbs_sel_i[3]
port 643 nsew
rlabel metal2 s 5234 -960 5346 480 4 wbs_stb_i
port 644 nsew
rlabel metal2 s 6430 -960 6542 480 4 wbs_we_i
port 645 nsew
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
