magic
tech sky130A
magscale 1 2
timestamp 1638581489
<< obsli1 >>
rect 1104 1377 141312 142001
<< obsm1 >>
rect 106 960 142310 142032
<< metal2 >>
rect 570 143820 626 144620
rect 1766 143820 1822 144620
rect 3054 143820 3110 144620
rect 4250 143820 4306 144620
rect 5538 143820 5594 144620
rect 6734 143820 6790 144620
rect 8022 143820 8078 144620
rect 9310 143820 9366 144620
rect 10506 143820 10562 144620
rect 11794 143820 11850 144620
rect 12990 143820 13046 144620
rect 14278 143820 14334 144620
rect 15566 143820 15622 144620
rect 16762 143820 16818 144620
rect 18050 143820 18106 144620
rect 19246 143820 19302 144620
rect 20534 143820 20590 144620
rect 21730 143820 21786 144620
rect 23018 143820 23074 144620
rect 24306 143820 24362 144620
rect 25502 143820 25558 144620
rect 26790 143820 26846 144620
rect 27986 143820 28042 144620
rect 29274 143820 29330 144620
rect 30562 143820 30618 144620
rect 31758 143820 31814 144620
rect 33046 143820 33102 144620
rect 34242 143820 34298 144620
rect 35530 143820 35586 144620
rect 36818 143820 36874 144620
rect 38014 143820 38070 144620
rect 39302 143820 39358 144620
rect 40498 143820 40554 144620
rect 41786 143820 41842 144620
rect 42982 143820 43038 144620
rect 44270 143820 44326 144620
rect 45558 143820 45614 144620
rect 46754 143820 46810 144620
rect 48042 143820 48098 144620
rect 49238 143820 49294 144620
rect 50526 143820 50582 144620
rect 51814 143820 51870 144620
rect 53010 143820 53066 144620
rect 54298 143820 54354 144620
rect 55494 143820 55550 144620
rect 56782 143820 56838 144620
rect 58070 143820 58126 144620
rect 59266 143820 59322 144620
rect 60554 143820 60610 144620
rect 61750 143820 61806 144620
rect 63038 143820 63094 144620
rect 64234 143820 64290 144620
rect 65522 143820 65578 144620
rect 66810 143820 66866 144620
rect 68006 143820 68062 144620
rect 69294 143820 69350 144620
rect 70490 143820 70546 144620
rect 71778 143820 71834 144620
rect 73066 143820 73122 144620
rect 74262 143820 74318 144620
rect 75550 143820 75606 144620
rect 76746 143820 76802 144620
rect 78034 143820 78090 144620
rect 79322 143820 79378 144620
rect 80518 143820 80574 144620
rect 81806 143820 81862 144620
rect 83002 143820 83058 144620
rect 84290 143820 84346 144620
rect 85486 143820 85542 144620
rect 86774 143820 86830 144620
rect 88062 143820 88118 144620
rect 89258 143820 89314 144620
rect 90546 143820 90602 144620
rect 91742 143820 91798 144620
rect 93030 143820 93086 144620
rect 94318 143820 94374 144620
rect 95514 143820 95570 144620
rect 96802 143820 96858 144620
rect 97998 143820 98054 144620
rect 99286 143820 99342 144620
rect 100574 143820 100630 144620
rect 101770 143820 101826 144620
rect 103058 143820 103114 144620
rect 104254 143820 104310 144620
rect 105542 143820 105598 144620
rect 106738 143820 106794 144620
rect 108026 143820 108082 144620
rect 109314 143820 109370 144620
rect 110510 143820 110566 144620
rect 111798 143820 111854 144620
rect 112994 143820 113050 144620
rect 114282 143820 114338 144620
rect 115570 143820 115626 144620
rect 116766 143820 116822 144620
rect 118054 143820 118110 144620
rect 119250 143820 119306 144620
rect 120538 143820 120594 144620
rect 121826 143820 121882 144620
rect 123022 143820 123078 144620
rect 124310 143820 124366 144620
rect 125506 143820 125562 144620
rect 126794 143820 126850 144620
rect 127990 143820 128046 144620
rect 129278 143820 129334 144620
rect 130566 143820 130622 144620
rect 131762 143820 131818 144620
rect 133050 143820 133106 144620
rect 134246 143820 134302 144620
rect 135534 143820 135590 144620
rect 136822 143820 136878 144620
rect 138018 143820 138074 144620
rect 139306 143820 139362 144620
rect 140502 143820 140558 144620
rect 141790 143820 141846 144620
rect 110 0 166 800
rect 386 0 442 800
rect 662 0 718 800
rect 938 0 994 800
rect 1214 0 1270 800
rect 1490 0 1546 800
rect 1766 0 1822 800
rect 2042 0 2098 800
rect 2410 0 2466 800
rect 2686 0 2742 800
rect 2962 0 3018 800
rect 3238 0 3294 800
rect 3514 0 3570 800
rect 3790 0 3846 800
rect 4066 0 4122 800
rect 4434 0 4490 800
rect 4710 0 4766 800
rect 4986 0 5042 800
rect 5262 0 5318 800
rect 5538 0 5594 800
rect 5814 0 5870 800
rect 6090 0 6146 800
rect 6458 0 6514 800
rect 6734 0 6790 800
rect 7010 0 7066 800
rect 7286 0 7342 800
rect 7562 0 7618 800
rect 7838 0 7894 800
rect 8114 0 8170 800
rect 8482 0 8538 800
rect 8758 0 8814 800
rect 9034 0 9090 800
rect 9310 0 9366 800
rect 9586 0 9642 800
rect 9862 0 9918 800
rect 10138 0 10194 800
rect 10506 0 10562 800
rect 10782 0 10838 800
rect 11058 0 11114 800
rect 11334 0 11390 800
rect 11610 0 11666 800
rect 11886 0 11942 800
rect 12162 0 12218 800
rect 12530 0 12586 800
rect 12806 0 12862 800
rect 13082 0 13138 800
rect 13358 0 13414 800
rect 13634 0 13690 800
rect 13910 0 13966 800
rect 14186 0 14242 800
rect 14554 0 14610 800
rect 14830 0 14886 800
rect 15106 0 15162 800
rect 15382 0 15438 800
rect 15658 0 15714 800
rect 15934 0 15990 800
rect 16210 0 16266 800
rect 16578 0 16634 800
rect 16854 0 16910 800
rect 17130 0 17186 800
rect 17406 0 17462 800
rect 17682 0 17738 800
rect 17958 0 18014 800
rect 18234 0 18290 800
rect 18602 0 18658 800
rect 18878 0 18934 800
rect 19154 0 19210 800
rect 19430 0 19486 800
rect 19706 0 19762 800
rect 19982 0 20038 800
rect 20258 0 20314 800
rect 20626 0 20682 800
rect 20902 0 20958 800
rect 21178 0 21234 800
rect 21454 0 21510 800
rect 21730 0 21786 800
rect 22006 0 22062 800
rect 22282 0 22338 800
rect 22650 0 22706 800
rect 22926 0 22982 800
rect 23202 0 23258 800
rect 23478 0 23534 800
rect 23754 0 23810 800
rect 24030 0 24086 800
rect 24306 0 24362 800
rect 24674 0 24730 800
rect 24950 0 25006 800
rect 25226 0 25282 800
rect 25502 0 25558 800
rect 25778 0 25834 800
rect 26054 0 26110 800
rect 26330 0 26386 800
rect 26698 0 26754 800
rect 26974 0 27030 800
rect 27250 0 27306 800
rect 27526 0 27582 800
rect 27802 0 27858 800
rect 28078 0 28134 800
rect 28354 0 28410 800
rect 28722 0 28778 800
rect 28998 0 29054 800
rect 29274 0 29330 800
rect 29550 0 29606 800
rect 29826 0 29882 800
rect 30102 0 30158 800
rect 30378 0 30434 800
rect 30746 0 30802 800
rect 31022 0 31078 800
rect 31298 0 31354 800
rect 31574 0 31630 800
rect 31850 0 31906 800
rect 32126 0 32182 800
rect 32402 0 32458 800
rect 32770 0 32826 800
rect 33046 0 33102 800
rect 33322 0 33378 800
rect 33598 0 33654 800
rect 33874 0 33930 800
rect 34150 0 34206 800
rect 34426 0 34482 800
rect 34794 0 34850 800
rect 35070 0 35126 800
rect 35346 0 35402 800
rect 35622 0 35678 800
rect 35898 0 35954 800
rect 36174 0 36230 800
rect 36450 0 36506 800
rect 36818 0 36874 800
rect 37094 0 37150 800
rect 37370 0 37426 800
rect 37646 0 37702 800
rect 37922 0 37978 800
rect 38198 0 38254 800
rect 38474 0 38530 800
rect 38842 0 38898 800
rect 39118 0 39174 800
rect 39394 0 39450 800
rect 39670 0 39726 800
rect 39946 0 40002 800
rect 40222 0 40278 800
rect 40498 0 40554 800
rect 40866 0 40922 800
rect 41142 0 41198 800
rect 41418 0 41474 800
rect 41694 0 41750 800
rect 41970 0 42026 800
rect 42246 0 42302 800
rect 42522 0 42578 800
rect 42890 0 42946 800
rect 43166 0 43222 800
rect 43442 0 43498 800
rect 43718 0 43774 800
rect 43994 0 44050 800
rect 44270 0 44326 800
rect 44546 0 44602 800
rect 44914 0 44970 800
rect 45190 0 45246 800
rect 45466 0 45522 800
rect 45742 0 45798 800
rect 46018 0 46074 800
rect 46294 0 46350 800
rect 46570 0 46626 800
rect 46938 0 46994 800
rect 47214 0 47270 800
rect 47490 0 47546 800
rect 47766 0 47822 800
rect 48042 0 48098 800
rect 48318 0 48374 800
rect 48594 0 48650 800
rect 48870 0 48926 800
rect 49238 0 49294 800
rect 49514 0 49570 800
rect 49790 0 49846 800
rect 50066 0 50122 800
rect 50342 0 50398 800
rect 50618 0 50674 800
rect 50894 0 50950 800
rect 51262 0 51318 800
rect 51538 0 51594 800
rect 51814 0 51870 800
rect 52090 0 52146 800
rect 52366 0 52422 800
rect 52642 0 52698 800
rect 52918 0 52974 800
rect 53286 0 53342 800
rect 53562 0 53618 800
rect 53838 0 53894 800
rect 54114 0 54170 800
rect 54390 0 54446 800
rect 54666 0 54722 800
rect 54942 0 54998 800
rect 55310 0 55366 800
rect 55586 0 55642 800
rect 55862 0 55918 800
rect 56138 0 56194 800
rect 56414 0 56470 800
rect 56690 0 56746 800
rect 56966 0 57022 800
rect 57334 0 57390 800
rect 57610 0 57666 800
rect 57886 0 57942 800
rect 58162 0 58218 800
rect 58438 0 58494 800
rect 58714 0 58770 800
rect 58990 0 59046 800
rect 59358 0 59414 800
rect 59634 0 59690 800
rect 59910 0 59966 800
rect 60186 0 60242 800
rect 60462 0 60518 800
rect 60738 0 60794 800
rect 61014 0 61070 800
rect 61382 0 61438 800
rect 61658 0 61714 800
rect 61934 0 61990 800
rect 62210 0 62266 800
rect 62486 0 62542 800
rect 62762 0 62818 800
rect 63038 0 63094 800
rect 63406 0 63462 800
rect 63682 0 63738 800
rect 63958 0 64014 800
rect 64234 0 64290 800
rect 64510 0 64566 800
rect 64786 0 64842 800
rect 65062 0 65118 800
rect 65430 0 65486 800
rect 65706 0 65762 800
rect 65982 0 66038 800
rect 66258 0 66314 800
rect 66534 0 66590 800
rect 66810 0 66866 800
rect 67086 0 67142 800
rect 67454 0 67510 800
rect 67730 0 67786 800
rect 68006 0 68062 800
rect 68282 0 68338 800
rect 68558 0 68614 800
rect 68834 0 68890 800
rect 69110 0 69166 800
rect 69478 0 69534 800
rect 69754 0 69810 800
rect 70030 0 70086 800
rect 70306 0 70362 800
rect 70582 0 70638 800
rect 70858 0 70914 800
rect 71134 0 71190 800
rect 71502 0 71558 800
rect 71778 0 71834 800
rect 72054 0 72110 800
rect 72330 0 72386 800
rect 72606 0 72662 800
rect 72882 0 72938 800
rect 73158 0 73214 800
rect 73526 0 73582 800
rect 73802 0 73858 800
rect 74078 0 74134 800
rect 74354 0 74410 800
rect 74630 0 74686 800
rect 74906 0 74962 800
rect 75182 0 75238 800
rect 75550 0 75606 800
rect 75826 0 75882 800
rect 76102 0 76158 800
rect 76378 0 76434 800
rect 76654 0 76710 800
rect 76930 0 76986 800
rect 77206 0 77262 800
rect 77574 0 77630 800
rect 77850 0 77906 800
rect 78126 0 78182 800
rect 78402 0 78458 800
rect 78678 0 78734 800
rect 78954 0 79010 800
rect 79230 0 79286 800
rect 79598 0 79654 800
rect 79874 0 79930 800
rect 80150 0 80206 800
rect 80426 0 80482 800
rect 80702 0 80758 800
rect 80978 0 81034 800
rect 81254 0 81310 800
rect 81622 0 81678 800
rect 81898 0 81954 800
rect 82174 0 82230 800
rect 82450 0 82506 800
rect 82726 0 82782 800
rect 83002 0 83058 800
rect 83278 0 83334 800
rect 83646 0 83702 800
rect 83922 0 83978 800
rect 84198 0 84254 800
rect 84474 0 84530 800
rect 84750 0 84806 800
rect 85026 0 85082 800
rect 85302 0 85358 800
rect 85670 0 85726 800
rect 85946 0 86002 800
rect 86222 0 86278 800
rect 86498 0 86554 800
rect 86774 0 86830 800
rect 87050 0 87106 800
rect 87326 0 87382 800
rect 87694 0 87750 800
rect 87970 0 88026 800
rect 88246 0 88302 800
rect 88522 0 88578 800
rect 88798 0 88854 800
rect 89074 0 89130 800
rect 89350 0 89406 800
rect 89718 0 89774 800
rect 89994 0 90050 800
rect 90270 0 90326 800
rect 90546 0 90602 800
rect 90822 0 90878 800
rect 91098 0 91154 800
rect 91374 0 91430 800
rect 91742 0 91798 800
rect 92018 0 92074 800
rect 92294 0 92350 800
rect 92570 0 92626 800
rect 92846 0 92902 800
rect 93122 0 93178 800
rect 93398 0 93454 800
rect 93766 0 93822 800
rect 94042 0 94098 800
rect 94318 0 94374 800
rect 94594 0 94650 800
rect 94870 0 94926 800
rect 95146 0 95202 800
rect 95422 0 95478 800
rect 95698 0 95754 800
rect 96066 0 96122 800
rect 96342 0 96398 800
rect 96618 0 96674 800
rect 96894 0 96950 800
rect 97170 0 97226 800
rect 97446 0 97502 800
rect 97722 0 97778 800
rect 98090 0 98146 800
rect 98366 0 98422 800
rect 98642 0 98698 800
rect 98918 0 98974 800
rect 99194 0 99250 800
rect 99470 0 99526 800
rect 99746 0 99802 800
rect 100114 0 100170 800
rect 100390 0 100446 800
rect 100666 0 100722 800
rect 100942 0 100998 800
rect 101218 0 101274 800
rect 101494 0 101550 800
rect 101770 0 101826 800
rect 102138 0 102194 800
rect 102414 0 102470 800
rect 102690 0 102746 800
rect 102966 0 103022 800
rect 103242 0 103298 800
rect 103518 0 103574 800
rect 103794 0 103850 800
rect 104162 0 104218 800
rect 104438 0 104494 800
rect 104714 0 104770 800
rect 104990 0 105046 800
rect 105266 0 105322 800
rect 105542 0 105598 800
rect 105818 0 105874 800
rect 106186 0 106242 800
rect 106462 0 106518 800
rect 106738 0 106794 800
rect 107014 0 107070 800
rect 107290 0 107346 800
rect 107566 0 107622 800
rect 107842 0 107898 800
rect 108210 0 108266 800
rect 108486 0 108542 800
rect 108762 0 108818 800
rect 109038 0 109094 800
rect 109314 0 109370 800
rect 109590 0 109646 800
rect 109866 0 109922 800
rect 110234 0 110290 800
rect 110510 0 110566 800
rect 110786 0 110842 800
rect 111062 0 111118 800
rect 111338 0 111394 800
rect 111614 0 111670 800
rect 111890 0 111946 800
rect 112258 0 112314 800
rect 112534 0 112590 800
rect 112810 0 112866 800
rect 113086 0 113142 800
rect 113362 0 113418 800
rect 113638 0 113694 800
rect 113914 0 113970 800
rect 114282 0 114338 800
rect 114558 0 114614 800
rect 114834 0 114890 800
rect 115110 0 115166 800
rect 115386 0 115442 800
rect 115662 0 115718 800
rect 115938 0 115994 800
rect 116306 0 116362 800
rect 116582 0 116638 800
rect 116858 0 116914 800
rect 117134 0 117190 800
rect 117410 0 117466 800
rect 117686 0 117742 800
rect 117962 0 118018 800
rect 118330 0 118386 800
rect 118606 0 118662 800
rect 118882 0 118938 800
rect 119158 0 119214 800
rect 119434 0 119490 800
rect 119710 0 119766 800
rect 119986 0 120042 800
rect 120354 0 120410 800
rect 120630 0 120686 800
rect 120906 0 120962 800
rect 121182 0 121238 800
rect 121458 0 121514 800
rect 121734 0 121790 800
rect 122010 0 122066 800
rect 122378 0 122434 800
rect 122654 0 122710 800
rect 122930 0 122986 800
rect 123206 0 123262 800
rect 123482 0 123538 800
rect 123758 0 123814 800
rect 124034 0 124090 800
rect 124402 0 124458 800
rect 124678 0 124734 800
rect 124954 0 125010 800
rect 125230 0 125286 800
rect 125506 0 125562 800
rect 125782 0 125838 800
rect 126058 0 126114 800
rect 126426 0 126482 800
rect 126702 0 126758 800
rect 126978 0 127034 800
rect 127254 0 127310 800
rect 127530 0 127586 800
rect 127806 0 127862 800
rect 128082 0 128138 800
rect 128450 0 128506 800
rect 128726 0 128782 800
rect 129002 0 129058 800
rect 129278 0 129334 800
rect 129554 0 129610 800
rect 129830 0 129886 800
rect 130106 0 130162 800
rect 130474 0 130530 800
rect 130750 0 130806 800
rect 131026 0 131082 800
rect 131302 0 131358 800
rect 131578 0 131634 800
rect 131854 0 131910 800
rect 132130 0 132186 800
rect 132498 0 132554 800
rect 132774 0 132830 800
rect 133050 0 133106 800
rect 133326 0 133382 800
rect 133602 0 133658 800
rect 133878 0 133934 800
rect 134154 0 134210 800
rect 134522 0 134578 800
rect 134798 0 134854 800
rect 135074 0 135130 800
rect 135350 0 135406 800
rect 135626 0 135682 800
rect 135902 0 135958 800
rect 136178 0 136234 800
rect 136546 0 136602 800
rect 136822 0 136878 800
rect 137098 0 137154 800
rect 137374 0 137430 800
rect 137650 0 137706 800
rect 137926 0 137982 800
rect 138202 0 138258 800
rect 138570 0 138626 800
rect 138846 0 138902 800
rect 139122 0 139178 800
rect 139398 0 139454 800
rect 139674 0 139730 800
rect 139950 0 140006 800
rect 140226 0 140282 800
rect 140594 0 140650 800
rect 140870 0 140926 800
rect 141146 0 141202 800
rect 141422 0 141478 800
rect 141698 0 141754 800
rect 141974 0 142030 800
rect 142250 0 142306 800
<< obsm2 >>
rect 112 143764 514 143834
rect 682 143764 1710 143834
rect 1878 143764 2998 143834
rect 3166 143764 4194 143834
rect 4362 143764 5482 143834
rect 5650 143764 6678 143834
rect 6846 143764 7966 143834
rect 8134 143764 9254 143834
rect 9422 143764 10450 143834
rect 10618 143764 11738 143834
rect 11906 143764 12934 143834
rect 13102 143764 14222 143834
rect 14390 143764 15510 143834
rect 15678 143764 16706 143834
rect 16874 143764 17994 143834
rect 18162 143764 19190 143834
rect 19358 143764 20478 143834
rect 20646 143764 21674 143834
rect 21842 143764 22962 143834
rect 23130 143764 24250 143834
rect 24418 143764 25446 143834
rect 25614 143764 26734 143834
rect 26902 143764 27930 143834
rect 28098 143764 29218 143834
rect 29386 143764 30506 143834
rect 30674 143764 31702 143834
rect 31870 143764 32990 143834
rect 33158 143764 34186 143834
rect 34354 143764 35474 143834
rect 35642 143764 36762 143834
rect 36930 143764 37958 143834
rect 38126 143764 39246 143834
rect 39414 143764 40442 143834
rect 40610 143764 41730 143834
rect 41898 143764 42926 143834
rect 43094 143764 44214 143834
rect 44382 143764 45502 143834
rect 45670 143764 46698 143834
rect 46866 143764 47986 143834
rect 48154 143764 49182 143834
rect 49350 143764 50470 143834
rect 50638 143764 51758 143834
rect 51926 143764 52954 143834
rect 53122 143764 54242 143834
rect 54410 143764 55438 143834
rect 55606 143764 56726 143834
rect 56894 143764 58014 143834
rect 58182 143764 59210 143834
rect 59378 143764 60498 143834
rect 60666 143764 61694 143834
rect 61862 143764 62982 143834
rect 63150 143764 64178 143834
rect 64346 143764 65466 143834
rect 65634 143764 66754 143834
rect 66922 143764 67950 143834
rect 68118 143764 69238 143834
rect 69406 143764 70434 143834
rect 70602 143764 71722 143834
rect 71890 143764 73010 143834
rect 73178 143764 74206 143834
rect 74374 143764 75494 143834
rect 75662 143764 76690 143834
rect 76858 143764 77978 143834
rect 78146 143764 79266 143834
rect 79434 143764 80462 143834
rect 80630 143764 81750 143834
rect 81918 143764 82946 143834
rect 83114 143764 84234 143834
rect 84402 143764 85430 143834
rect 85598 143764 86718 143834
rect 86886 143764 88006 143834
rect 88174 143764 89202 143834
rect 89370 143764 90490 143834
rect 90658 143764 91686 143834
rect 91854 143764 92974 143834
rect 93142 143764 94262 143834
rect 94430 143764 95458 143834
rect 95626 143764 96746 143834
rect 96914 143764 97942 143834
rect 98110 143764 99230 143834
rect 99398 143764 100518 143834
rect 100686 143764 101714 143834
rect 101882 143764 103002 143834
rect 103170 143764 104198 143834
rect 104366 143764 105486 143834
rect 105654 143764 106682 143834
rect 106850 143764 107970 143834
rect 108138 143764 109258 143834
rect 109426 143764 110454 143834
rect 110622 143764 111742 143834
rect 111910 143764 112938 143834
rect 113106 143764 114226 143834
rect 114394 143764 115514 143834
rect 115682 143764 116710 143834
rect 116878 143764 117998 143834
rect 118166 143764 119194 143834
rect 119362 143764 120482 143834
rect 120650 143764 121770 143834
rect 121938 143764 122966 143834
rect 123134 143764 124254 143834
rect 124422 143764 125450 143834
rect 125618 143764 126738 143834
rect 126906 143764 127934 143834
rect 128102 143764 129222 143834
rect 129390 143764 130510 143834
rect 130678 143764 131706 143834
rect 131874 143764 132994 143834
rect 133162 143764 134190 143834
rect 134358 143764 135478 143834
rect 135646 143764 136766 143834
rect 136934 143764 137962 143834
rect 138130 143764 139250 143834
rect 139418 143764 140446 143834
rect 140614 143764 141734 143834
rect 141902 143764 142304 143834
rect 112 856 142304 143764
rect 222 734 330 856
rect 498 734 606 856
rect 774 734 882 856
rect 1050 734 1158 856
rect 1326 734 1434 856
rect 1602 734 1710 856
rect 1878 734 1986 856
rect 2154 734 2354 856
rect 2522 734 2630 856
rect 2798 734 2906 856
rect 3074 734 3182 856
rect 3350 734 3458 856
rect 3626 734 3734 856
rect 3902 734 4010 856
rect 4178 734 4378 856
rect 4546 734 4654 856
rect 4822 734 4930 856
rect 5098 734 5206 856
rect 5374 734 5482 856
rect 5650 734 5758 856
rect 5926 734 6034 856
rect 6202 734 6402 856
rect 6570 734 6678 856
rect 6846 734 6954 856
rect 7122 734 7230 856
rect 7398 734 7506 856
rect 7674 734 7782 856
rect 7950 734 8058 856
rect 8226 734 8426 856
rect 8594 734 8702 856
rect 8870 734 8978 856
rect 9146 734 9254 856
rect 9422 734 9530 856
rect 9698 734 9806 856
rect 9974 734 10082 856
rect 10250 734 10450 856
rect 10618 734 10726 856
rect 10894 734 11002 856
rect 11170 734 11278 856
rect 11446 734 11554 856
rect 11722 734 11830 856
rect 11998 734 12106 856
rect 12274 734 12474 856
rect 12642 734 12750 856
rect 12918 734 13026 856
rect 13194 734 13302 856
rect 13470 734 13578 856
rect 13746 734 13854 856
rect 14022 734 14130 856
rect 14298 734 14498 856
rect 14666 734 14774 856
rect 14942 734 15050 856
rect 15218 734 15326 856
rect 15494 734 15602 856
rect 15770 734 15878 856
rect 16046 734 16154 856
rect 16322 734 16522 856
rect 16690 734 16798 856
rect 16966 734 17074 856
rect 17242 734 17350 856
rect 17518 734 17626 856
rect 17794 734 17902 856
rect 18070 734 18178 856
rect 18346 734 18546 856
rect 18714 734 18822 856
rect 18990 734 19098 856
rect 19266 734 19374 856
rect 19542 734 19650 856
rect 19818 734 19926 856
rect 20094 734 20202 856
rect 20370 734 20570 856
rect 20738 734 20846 856
rect 21014 734 21122 856
rect 21290 734 21398 856
rect 21566 734 21674 856
rect 21842 734 21950 856
rect 22118 734 22226 856
rect 22394 734 22594 856
rect 22762 734 22870 856
rect 23038 734 23146 856
rect 23314 734 23422 856
rect 23590 734 23698 856
rect 23866 734 23974 856
rect 24142 734 24250 856
rect 24418 734 24618 856
rect 24786 734 24894 856
rect 25062 734 25170 856
rect 25338 734 25446 856
rect 25614 734 25722 856
rect 25890 734 25998 856
rect 26166 734 26274 856
rect 26442 734 26642 856
rect 26810 734 26918 856
rect 27086 734 27194 856
rect 27362 734 27470 856
rect 27638 734 27746 856
rect 27914 734 28022 856
rect 28190 734 28298 856
rect 28466 734 28666 856
rect 28834 734 28942 856
rect 29110 734 29218 856
rect 29386 734 29494 856
rect 29662 734 29770 856
rect 29938 734 30046 856
rect 30214 734 30322 856
rect 30490 734 30690 856
rect 30858 734 30966 856
rect 31134 734 31242 856
rect 31410 734 31518 856
rect 31686 734 31794 856
rect 31962 734 32070 856
rect 32238 734 32346 856
rect 32514 734 32714 856
rect 32882 734 32990 856
rect 33158 734 33266 856
rect 33434 734 33542 856
rect 33710 734 33818 856
rect 33986 734 34094 856
rect 34262 734 34370 856
rect 34538 734 34738 856
rect 34906 734 35014 856
rect 35182 734 35290 856
rect 35458 734 35566 856
rect 35734 734 35842 856
rect 36010 734 36118 856
rect 36286 734 36394 856
rect 36562 734 36762 856
rect 36930 734 37038 856
rect 37206 734 37314 856
rect 37482 734 37590 856
rect 37758 734 37866 856
rect 38034 734 38142 856
rect 38310 734 38418 856
rect 38586 734 38786 856
rect 38954 734 39062 856
rect 39230 734 39338 856
rect 39506 734 39614 856
rect 39782 734 39890 856
rect 40058 734 40166 856
rect 40334 734 40442 856
rect 40610 734 40810 856
rect 40978 734 41086 856
rect 41254 734 41362 856
rect 41530 734 41638 856
rect 41806 734 41914 856
rect 42082 734 42190 856
rect 42358 734 42466 856
rect 42634 734 42834 856
rect 43002 734 43110 856
rect 43278 734 43386 856
rect 43554 734 43662 856
rect 43830 734 43938 856
rect 44106 734 44214 856
rect 44382 734 44490 856
rect 44658 734 44858 856
rect 45026 734 45134 856
rect 45302 734 45410 856
rect 45578 734 45686 856
rect 45854 734 45962 856
rect 46130 734 46238 856
rect 46406 734 46514 856
rect 46682 734 46882 856
rect 47050 734 47158 856
rect 47326 734 47434 856
rect 47602 734 47710 856
rect 47878 734 47986 856
rect 48154 734 48262 856
rect 48430 734 48538 856
rect 48706 734 48814 856
rect 48982 734 49182 856
rect 49350 734 49458 856
rect 49626 734 49734 856
rect 49902 734 50010 856
rect 50178 734 50286 856
rect 50454 734 50562 856
rect 50730 734 50838 856
rect 51006 734 51206 856
rect 51374 734 51482 856
rect 51650 734 51758 856
rect 51926 734 52034 856
rect 52202 734 52310 856
rect 52478 734 52586 856
rect 52754 734 52862 856
rect 53030 734 53230 856
rect 53398 734 53506 856
rect 53674 734 53782 856
rect 53950 734 54058 856
rect 54226 734 54334 856
rect 54502 734 54610 856
rect 54778 734 54886 856
rect 55054 734 55254 856
rect 55422 734 55530 856
rect 55698 734 55806 856
rect 55974 734 56082 856
rect 56250 734 56358 856
rect 56526 734 56634 856
rect 56802 734 56910 856
rect 57078 734 57278 856
rect 57446 734 57554 856
rect 57722 734 57830 856
rect 57998 734 58106 856
rect 58274 734 58382 856
rect 58550 734 58658 856
rect 58826 734 58934 856
rect 59102 734 59302 856
rect 59470 734 59578 856
rect 59746 734 59854 856
rect 60022 734 60130 856
rect 60298 734 60406 856
rect 60574 734 60682 856
rect 60850 734 60958 856
rect 61126 734 61326 856
rect 61494 734 61602 856
rect 61770 734 61878 856
rect 62046 734 62154 856
rect 62322 734 62430 856
rect 62598 734 62706 856
rect 62874 734 62982 856
rect 63150 734 63350 856
rect 63518 734 63626 856
rect 63794 734 63902 856
rect 64070 734 64178 856
rect 64346 734 64454 856
rect 64622 734 64730 856
rect 64898 734 65006 856
rect 65174 734 65374 856
rect 65542 734 65650 856
rect 65818 734 65926 856
rect 66094 734 66202 856
rect 66370 734 66478 856
rect 66646 734 66754 856
rect 66922 734 67030 856
rect 67198 734 67398 856
rect 67566 734 67674 856
rect 67842 734 67950 856
rect 68118 734 68226 856
rect 68394 734 68502 856
rect 68670 734 68778 856
rect 68946 734 69054 856
rect 69222 734 69422 856
rect 69590 734 69698 856
rect 69866 734 69974 856
rect 70142 734 70250 856
rect 70418 734 70526 856
rect 70694 734 70802 856
rect 70970 734 71078 856
rect 71246 734 71446 856
rect 71614 734 71722 856
rect 71890 734 71998 856
rect 72166 734 72274 856
rect 72442 734 72550 856
rect 72718 734 72826 856
rect 72994 734 73102 856
rect 73270 734 73470 856
rect 73638 734 73746 856
rect 73914 734 74022 856
rect 74190 734 74298 856
rect 74466 734 74574 856
rect 74742 734 74850 856
rect 75018 734 75126 856
rect 75294 734 75494 856
rect 75662 734 75770 856
rect 75938 734 76046 856
rect 76214 734 76322 856
rect 76490 734 76598 856
rect 76766 734 76874 856
rect 77042 734 77150 856
rect 77318 734 77518 856
rect 77686 734 77794 856
rect 77962 734 78070 856
rect 78238 734 78346 856
rect 78514 734 78622 856
rect 78790 734 78898 856
rect 79066 734 79174 856
rect 79342 734 79542 856
rect 79710 734 79818 856
rect 79986 734 80094 856
rect 80262 734 80370 856
rect 80538 734 80646 856
rect 80814 734 80922 856
rect 81090 734 81198 856
rect 81366 734 81566 856
rect 81734 734 81842 856
rect 82010 734 82118 856
rect 82286 734 82394 856
rect 82562 734 82670 856
rect 82838 734 82946 856
rect 83114 734 83222 856
rect 83390 734 83590 856
rect 83758 734 83866 856
rect 84034 734 84142 856
rect 84310 734 84418 856
rect 84586 734 84694 856
rect 84862 734 84970 856
rect 85138 734 85246 856
rect 85414 734 85614 856
rect 85782 734 85890 856
rect 86058 734 86166 856
rect 86334 734 86442 856
rect 86610 734 86718 856
rect 86886 734 86994 856
rect 87162 734 87270 856
rect 87438 734 87638 856
rect 87806 734 87914 856
rect 88082 734 88190 856
rect 88358 734 88466 856
rect 88634 734 88742 856
rect 88910 734 89018 856
rect 89186 734 89294 856
rect 89462 734 89662 856
rect 89830 734 89938 856
rect 90106 734 90214 856
rect 90382 734 90490 856
rect 90658 734 90766 856
rect 90934 734 91042 856
rect 91210 734 91318 856
rect 91486 734 91686 856
rect 91854 734 91962 856
rect 92130 734 92238 856
rect 92406 734 92514 856
rect 92682 734 92790 856
rect 92958 734 93066 856
rect 93234 734 93342 856
rect 93510 734 93710 856
rect 93878 734 93986 856
rect 94154 734 94262 856
rect 94430 734 94538 856
rect 94706 734 94814 856
rect 94982 734 95090 856
rect 95258 734 95366 856
rect 95534 734 95642 856
rect 95810 734 96010 856
rect 96178 734 96286 856
rect 96454 734 96562 856
rect 96730 734 96838 856
rect 97006 734 97114 856
rect 97282 734 97390 856
rect 97558 734 97666 856
rect 97834 734 98034 856
rect 98202 734 98310 856
rect 98478 734 98586 856
rect 98754 734 98862 856
rect 99030 734 99138 856
rect 99306 734 99414 856
rect 99582 734 99690 856
rect 99858 734 100058 856
rect 100226 734 100334 856
rect 100502 734 100610 856
rect 100778 734 100886 856
rect 101054 734 101162 856
rect 101330 734 101438 856
rect 101606 734 101714 856
rect 101882 734 102082 856
rect 102250 734 102358 856
rect 102526 734 102634 856
rect 102802 734 102910 856
rect 103078 734 103186 856
rect 103354 734 103462 856
rect 103630 734 103738 856
rect 103906 734 104106 856
rect 104274 734 104382 856
rect 104550 734 104658 856
rect 104826 734 104934 856
rect 105102 734 105210 856
rect 105378 734 105486 856
rect 105654 734 105762 856
rect 105930 734 106130 856
rect 106298 734 106406 856
rect 106574 734 106682 856
rect 106850 734 106958 856
rect 107126 734 107234 856
rect 107402 734 107510 856
rect 107678 734 107786 856
rect 107954 734 108154 856
rect 108322 734 108430 856
rect 108598 734 108706 856
rect 108874 734 108982 856
rect 109150 734 109258 856
rect 109426 734 109534 856
rect 109702 734 109810 856
rect 109978 734 110178 856
rect 110346 734 110454 856
rect 110622 734 110730 856
rect 110898 734 111006 856
rect 111174 734 111282 856
rect 111450 734 111558 856
rect 111726 734 111834 856
rect 112002 734 112202 856
rect 112370 734 112478 856
rect 112646 734 112754 856
rect 112922 734 113030 856
rect 113198 734 113306 856
rect 113474 734 113582 856
rect 113750 734 113858 856
rect 114026 734 114226 856
rect 114394 734 114502 856
rect 114670 734 114778 856
rect 114946 734 115054 856
rect 115222 734 115330 856
rect 115498 734 115606 856
rect 115774 734 115882 856
rect 116050 734 116250 856
rect 116418 734 116526 856
rect 116694 734 116802 856
rect 116970 734 117078 856
rect 117246 734 117354 856
rect 117522 734 117630 856
rect 117798 734 117906 856
rect 118074 734 118274 856
rect 118442 734 118550 856
rect 118718 734 118826 856
rect 118994 734 119102 856
rect 119270 734 119378 856
rect 119546 734 119654 856
rect 119822 734 119930 856
rect 120098 734 120298 856
rect 120466 734 120574 856
rect 120742 734 120850 856
rect 121018 734 121126 856
rect 121294 734 121402 856
rect 121570 734 121678 856
rect 121846 734 121954 856
rect 122122 734 122322 856
rect 122490 734 122598 856
rect 122766 734 122874 856
rect 123042 734 123150 856
rect 123318 734 123426 856
rect 123594 734 123702 856
rect 123870 734 123978 856
rect 124146 734 124346 856
rect 124514 734 124622 856
rect 124790 734 124898 856
rect 125066 734 125174 856
rect 125342 734 125450 856
rect 125618 734 125726 856
rect 125894 734 126002 856
rect 126170 734 126370 856
rect 126538 734 126646 856
rect 126814 734 126922 856
rect 127090 734 127198 856
rect 127366 734 127474 856
rect 127642 734 127750 856
rect 127918 734 128026 856
rect 128194 734 128394 856
rect 128562 734 128670 856
rect 128838 734 128946 856
rect 129114 734 129222 856
rect 129390 734 129498 856
rect 129666 734 129774 856
rect 129942 734 130050 856
rect 130218 734 130418 856
rect 130586 734 130694 856
rect 130862 734 130970 856
rect 131138 734 131246 856
rect 131414 734 131522 856
rect 131690 734 131798 856
rect 131966 734 132074 856
rect 132242 734 132442 856
rect 132610 734 132718 856
rect 132886 734 132994 856
rect 133162 734 133270 856
rect 133438 734 133546 856
rect 133714 734 133822 856
rect 133990 734 134098 856
rect 134266 734 134466 856
rect 134634 734 134742 856
rect 134910 734 135018 856
rect 135186 734 135294 856
rect 135462 734 135570 856
rect 135738 734 135846 856
rect 136014 734 136122 856
rect 136290 734 136490 856
rect 136658 734 136766 856
rect 136934 734 137042 856
rect 137210 734 137318 856
rect 137486 734 137594 856
rect 137762 734 137870 856
rect 138038 734 138146 856
rect 138314 734 138514 856
rect 138682 734 138790 856
rect 138958 734 139066 856
rect 139234 734 139342 856
rect 139510 734 139618 856
rect 139786 734 139894 856
rect 140062 734 140170 856
rect 140338 734 140538 856
rect 140706 734 140814 856
rect 140982 734 141090 856
rect 141258 734 141366 856
rect 141534 734 141642 856
rect 141810 734 141918 856
rect 142086 734 142194 856
<< obsm3 >>
rect 1485 1803 140379 142017
<< metal4 >>
rect 4208 2128 4528 142032
rect 19568 2128 19888 142032
rect 34928 2128 35248 142032
rect 50288 2128 50608 142032
rect 65648 2128 65968 142032
rect 81008 2128 81328 142032
rect 96368 2128 96688 142032
rect 111728 2128 112048 142032
rect 127088 2128 127408 142032
<< obsm4 >>
rect 4843 2619 19488 130253
rect 19968 2619 34848 130253
rect 35328 2619 50208 130253
rect 50688 2619 65568 130253
rect 66048 2619 80928 130253
rect 81408 2619 96288 130253
rect 96768 2619 111648 130253
rect 112128 2619 127008 130253
rect 127488 2619 131133 130253
<< labels >>
rlabel metal2 s 570 143820 626 144620 6 io_in[0]
port 1 nsew signal input
rlabel metal2 s 38014 143820 38070 144620 6 io_in[10]
port 2 nsew signal input
rlabel metal2 s 41786 143820 41842 144620 6 io_in[11]
port 3 nsew signal input
rlabel metal2 s 45558 143820 45614 144620 6 io_in[12]
port 4 nsew signal input
rlabel metal2 s 49238 143820 49294 144620 6 io_in[13]
port 5 nsew signal input
rlabel metal2 s 53010 143820 53066 144620 6 io_in[14]
port 6 nsew signal input
rlabel metal2 s 56782 143820 56838 144620 6 io_in[15]
port 7 nsew signal input
rlabel metal2 s 60554 143820 60610 144620 6 io_in[16]
port 8 nsew signal input
rlabel metal2 s 64234 143820 64290 144620 6 io_in[17]
port 9 nsew signal input
rlabel metal2 s 68006 143820 68062 144620 6 io_in[18]
port 10 nsew signal input
rlabel metal2 s 71778 143820 71834 144620 6 io_in[19]
port 11 nsew signal input
rlabel metal2 s 4250 143820 4306 144620 6 io_in[1]
port 12 nsew signal input
rlabel metal2 s 75550 143820 75606 144620 6 io_in[20]
port 13 nsew signal input
rlabel metal2 s 79322 143820 79378 144620 6 io_in[21]
port 14 nsew signal input
rlabel metal2 s 83002 143820 83058 144620 6 io_in[22]
port 15 nsew signal input
rlabel metal2 s 86774 143820 86830 144620 6 io_in[23]
port 16 nsew signal input
rlabel metal2 s 90546 143820 90602 144620 6 io_in[24]
port 17 nsew signal input
rlabel metal2 s 94318 143820 94374 144620 6 io_in[25]
port 18 nsew signal input
rlabel metal2 s 97998 143820 98054 144620 6 io_in[26]
port 19 nsew signal input
rlabel metal2 s 101770 143820 101826 144620 6 io_in[27]
port 20 nsew signal input
rlabel metal2 s 105542 143820 105598 144620 6 io_in[28]
port 21 nsew signal input
rlabel metal2 s 109314 143820 109370 144620 6 io_in[29]
port 22 nsew signal input
rlabel metal2 s 8022 143820 8078 144620 6 io_in[2]
port 23 nsew signal input
rlabel metal2 s 112994 143820 113050 144620 6 io_in[30]
port 24 nsew signal input
rlabel metal2 s 116766 143820 116822 144620 6 io_in[31]
port 25 nsew signal input
rlabel metal2 s 120538 143820 120594 144620 6 io_in[32]
port 26 nsew signal input
rlabel metal2 s 124310 143820 124366 144620 6 io_in[33]
port 27 nsew signal input
rlabel metal2 s 127990 143820 128046 144620 6 io_in[34]
port 28 nsew signal input
rlabel metal2 s 131762 143820 131818 144620 6 io_in[35]
port 29 nsew signal input
rlabel metal2 s 135534 143820 135590 144620 6 io_in[36]
port 30 nsew signal input
rlabel metal2 s 139306 143820 139362 144620 6 io_in[37]
port 31 nsew signal input
rlabel metal2 s 11794 143820 11850 144620 6 io_in[3]
port 32 nsew signal input
rlabel metal2 s 15566 143820 15622 144620 6 io_in[4]
port 33 nsew signal input
rlabel metal2 s 19246 143820 19302 144620 6 io_in[5]
port 34 nsew signal input
rlabel metal2 s 23018 143820 23074 144620 6 io_in[6]
port 35 nsew signal input
rlabel metal2 s 26790 143820 26846 144620 6 io_in[7]
port 36 nsew signal input
rlabel metal2 s 30562 143820 30618 144620 6 io_in[8]
port 37 nsew signal input
rlabel metal2 s 34242 143820 34298 144620 6 io_in[9]
port 38 nsew signal input
rlabel metal2 s 1766 143820 1822 144620 6 io_oeb[0]
port 39 nsew signal output
rlabel metal2 s 39302 143820 39358 144620 6 io_oeb[10]
port 40 nsew signal output
rlabel metal2 s 42982 143820 43038 144620 6 io_oeb[11]
port 41 nsew signal output
rlabel metal2 s 46754 143820 46810 144620 6 io_oeb[12]
port 42 nsew signal output
rlabel metal2 s 50526 143820 50582 144620 6 io_oeb[13]
port 43 nsew signal output
rlabel metal2 s 54298 143820 54354 144620 6 io_oeb[14]
port 44 nsew signal output
rlabel metal2 s 58070 143820 58126 144620 6 io_oeb[15]
port 45 nsew signal output
rlabel metal2 s 61750 143820 61806 144620 6 io_oeb[16]
port 46 nsew signal output
rlabel metal2 s 65522 143820 65578 144620 6 io_oeb[17]
port 47 nsew signal output
rlabel metal2 s 69294 143820 69350 144620 6 io_oeb[18]
port 48 nsew signal output
rlabel metal2 s 73066 143820 73122 144620 6 io_oeb[19]
port 49 nsew signal output
rlabel metal2 s 5538 143820 5594 144620 6 io_oeb[1]
port 50 nsew signal output
rlabel metal2 s 76746 143820 76802 144620 6 io_oeb[20]
port 51 nsew signal output
rlabel metal2 s 80518 143820 80574 144620 6 io_oeb[21]
port 52 nsew signal output
rlabel metal2 s 84290 143820 84346 144620 6 io_oeb[22]
port 53 nsew signal output
rlabel metal2 s 88062 143820 88118 144620 6 io_oeb[23]
port 54 nsew signal output
rlabel metal2 s 91742 143820 91798 144620 6 io_oeb[24]
port 55 nsew signal output
rlabel metal2 s 95514 143820 95570 144620 6 io_oeb[25]
port 56 nsew signal output
rlabel metal2 s 99286 143820 99342 144620 6 io_oeb[26]
port 57 nsew signal output
rlabel metal2 s 103058 143820 103114 144620 6 io_oeb[27]
port 58 nsew signal output
rlabel metal2 s 106738 143820 106794 144620 6 io_oeb[28]
port 59 nsew signal output
rlabel metal2 s 110510 143820 110566 144620 6 io_oeb[29]
port 60 nsew signal output
rlabel metal2 s 9310 143820 9366 144620 6 io_oeb[2]
port 61 nsew signal output
rlabel metal2 s 114282 143820 114338 144620 6 io_oeb[30]
port 62 nsew signal output
rlabel metal2 s 118054 143820 118110 144620 6 io_oeb[31]
port 63 nsew signal output
rlabel metal2 s 121826 143820 121882 144620 6 io_oeb[32]
port 64 nsew signal output
rlabel metal2 s 125506 143820 125562 144620 6 io_oeb[33]
port 65 nsew signal output
rlabel metal2 s 129278 143820 129334 144620 6 io_oeb[34]
port 66 nsew signal output
rlabel metal2 s 133050 143820 133106 144620 6 io_oeb[35]
port 67 nsew signal output
rlabel metal2 s 136822 143820 136878 144620 6 io_oeb[36]
port 68 nsew signal output
rlabel metal2 s 140502 143820 140558 144620 6 io_oeb[37]
port 69 nsew signal output
rlabel metal2 s 12990 143820 13046 144620 6 io_oeb[3]
port 70 nsew signal output
rlabel metal2 s 16762 143820 16818 144620 6 io_oeb[4]
port 71 nsew signal output
rlabel metal2 s 20534 143820 20590 144620 6 io_oeb[5]
port 72 nsew signal output
rlabel metal2 s 24306 143820 24362 144620 6 io_oeb[6]
port 73 nsew signal output
rlabel metal2 s 27986 143820 28042 144620 6 io_oeb[7]
port 74 nsew signal output
rlabel metal2 s 31758 143820 31814 144620 6 io_oeb[8]
port 75 nsew signal output
rlabel metal2 s 35530 143820 35586 144620 6 io_oeb[9]
port 76 nsew signal output
rlabel metal2 s 3054 143820 3110 144620 6 io_out[0]
port 77 nsew signal output
rlabel metal2 s 40498 143820 40554 144620 6 io_out[10]
port 78 nsew signal output
rlabel metal2 s 44270 143820 44326 144620 6 io_out[11]
port 79 nsew signal output
rlabel metal2 s 48042 143820 48098 144620 6 io_out[12]
port 80 nsew signal output
rlabel metal2 s 51814 143820 51870 144620 6 io_out[13]
port 81 nsew signal output
rlabel metal2 s 55494 143820 55550 144620 6 io_out[14]
port 82 nsew signal output
rlabel metal2 s 59266 143820 59322 144620 6 io_out[15]
port 83 nsew signal output
rlabel metal2 s 63038 143820 63094 144620 6 io_out[16]
port 84 nsew signal output
rlabel metal2 s 66810 143820 66866 144620 6 io_out[17]
port 85 nsew signal output
rlabel metal2 s 70490 143820 70546 144620 6 io_out[18]
port 86 nsew signal output
rlabel metal2 s 74262 143820 74318 144620 6 io_out[19]
port 87 nsew signal output
rlabel metal2 s 6734 143820 6790 144620 6 io_out[1]
port 88 nsew signal output
rlabel metal2 s 78034 143820 78090 144620 6 io_out[20]
port 89 nsew signal output
rlabel metal2 s 81806 143820 81862 144620 6 io_out[21]
port 90 nsew signal output
rlabel metal2 s 85486 143820 85542 144620 6 io_out[22]
port 91 nsew signal output
rlabel metal2 s 89258 143820 89314 144620 6 io_out[23]
port 92 nsew signal output
rlabel metal2 s 93030 143820 93086 144620 6 io_out[24]
port 93 nsew signal output
rlabel metal2 s 96802 143820 96858 144620 6 io_out[25]
port 94 nsew signal output
rlabel metal2 s 100574 143820 100630 144620 6 io_out[26]
port 95 nsew signal output
rlabel metal2 s 104254 143820 104310 144620 6 io_out[27]
port 96 nsew signal output
rlabel metal2 s 108026 143820 108082 144620 6 io_out[28]
port 97 nsew signal output
rlabel metal2 s 111798 143820 111854 144620 6 io_out[29]
port 98 nsew signal output
rlabel metal2 s 10506 143820 10562 144620 6 io_out[2]
port 99 nsew signal output
rlabel metal2 s 115570 143820 115626 144620 6 io_out[30]
port 100 nsew signal output
rlabel metal2 s 119250 143820 119306 144620 6 io_out[31]
port 101 nsew signal output
rlabel metal2 s 123022 143820 123078 144620 6 io_out[32]
port 102 nsew signal output
rlabel metal2 s 126794 143820 126850 144620 6 io_out[33]
port 103 nsew signal output
rlabel metal2 s 130566 143820 130622 144620 6 io_out[34]
port 104 nsew signal output
rlabel metal2 s 134246 143820 134302 144620 6 io_out[35]
port 105 nsew signal output
rlabel metal2 s 138018 143820 138074 144620 6 io_out[36]
port 106 nsew signal output
rlabel metal2 s 141790 143820 141846 144620 6 io_out[37]
port 107 nsew signal output
rlabel metal2 s 14278 143820 14334 144620 6 io_out[3]
port 108 nsew signal output
rlabel metal2 s 18050 143820 18106 144620 6 io_out[4]
port 109 nsew signal output
rlabel metal2 s 21730 143820 21786 144620 6 io_out[5]
port 110 nsew signal output
rlabel metal2 s 25502 143820 25558 144620 6 io_out[6]
port 111 nsew signal output
rlabel metal2 s 29274 143820 29330 144620 6 io_out[7]
port 112 nsew signal output
rlabel metal2 s 33046 143820 33102 144620 6 io_out[8]
port 113 nsew signal output
rlabel metal2 s 36818 143820 36874 144620 6 io_out[9]
port 114 nsew signal output
rlabel metal2 s 141698 0 141754 800 6 irq[0]
port 115 nsew signal output
rlabel metal2 s 141974 0 142030 800 6 irq[1]
port 116 nsew signal output
rlabel metal2 s 142250 0 142306 800 6 irq[2]
port 117 nsew signal output
rlabel metal2 s 30746 0 30802 800 6 la_data_in[0]
port 118 nsew signal input
rlabel metal2 s 117410 0 117466 800 6 la_data_in[100]
port 119 nsew signal input
rlabel metal2 s 118330 0 118386 800 6 la_data_in[101]
port 120 nsew signal input
rlabel metal2 s 119158 0 119214 800 6 la_data_in[102]
port 121 nsew signal input
rlabel metal2 s 119986 0 120042 800 6 la_data_in[103]
port 122 nsew signal input
rlabel metal2 s 120906 0 120962 800 6 la_data_in[104]
port 123 nsew signal input
rlabel metal2 s 121734 0 121790 800 6 la_data_in[105]
port 124 nsew signal input
rlabel metal2 s 122654 0 122710 800 6 la_data_in[106]
port 125 nsew signal input
rlabel metal2 s 123482 0 123538 800 6 la_data_in[107]
port 126 nsew signal input
rlabel metal2 s 124402 0 124458 800 6 la_data_in[108]
port 127 nsew signal input
rlabel metal2 s 125230 0 125286 800 6 la_data_in[109]
port 128 nsew signal input
rlabel metal2 s 39394 0 39450 800 6 la_data_in[10]
port 129 nsew signal input
rlabel metal2 s 126058 0 126114 800 6 la_data_in[110]
port 130 nsew signal input
rlabel metal2 s 126978 0 127034 800 6 la_data_in[111]
port 131 nsew signal input
rlabel metal2 s 127806 0 127862 800 6 la_data_in[112]
port 132 nsew signal input
rlabel metal2 s 128726 0 128782 800 6 la_data_in[113]
port 133 nsew signal input
rlabel metal2 s 129554 0 129610 800 6 la_data_in[114]
port 134 nsew signal input
rlabel metal2 s 130474 0 130530 800 6 la_data_in[115]
port 135 nsew signal input
rlabel metal2 s 131302 0 131358 800 6 la_data_in[116]
port 136 nsew signal input
rlabel metal2 s 132130 0 132186 800 6 la_data_in[117]
port 137 nsew signal input
rlabel metal2 s 133050 0 133106 800 6 la_data_in[118]
port 138 nsew signal input
rlabel metal2 s 133878 0 133934 800 6 la_data_in[119]
port 139 nsew signal input
rlabel metal2 s 40222 0 40278 800 6 la_data_in[11]
port 140 nsew signal input
rlabel metal2 s 134798 0 134854 800 6 la_data_in[120]
port 141 nsew signal input
rlabel metal2 s 135626 0 135682 800 6 la_data_in[121]
port 142 nsew signal input
rlabel metal2 s 136546 0 136602 800 6 la_data_in[122]
port 143 nsew signal input
rlabel metal2 s 137374 0 137430 800 6 la_data_in[123]
port 144 nsew signal input
rlabel metal2 s 138202 0 138258 800 6 la_data_in[124]
port 145 nsew signal input
rlabel metal2 s 139122 0 139178 800 6 la_data_in[125]
port 146 nsew signal input
rlabel metal2 s 139950 0 140006 800 6 la_data_in[126]
port 147 nsew signal input
rlabel metal2 s 140870 0 140926 800 6 la_data_in[127]
port 148 nsew signal input
rlabel metal2 s 41142 0 41198 800 6 la_data_in[12]
port 149 nsew signal input
rlabel metal2 s 41970 0 42026 800 6 la_data_in[13]
port 150 nsew signal input
rlabel metal2 s 42890 0 42946 800 6 la_data_in[14]
port 151 nsew signal input
rlabel metal2 s 43718 0 43774 800 6 la_data_in[15]
port 152 nsew signal input
rlabel metal2 s 44546 0 44602 800 6 la_data_in[16]
port 153 nsew signal input
rlabel metal2 s 45466 0 45522 800 6 la_data_in[17]
port 154 nsew signal input
rlabel metal2 s 46294 0 46350 800 6 la_data_in[18]
port 155 nsew signal input
rlabel metal2 s 47214 0 47270 800 6 la_data_in[19]
port 156 nsew signal input
rlabel metal2 s 31574 0 31630 800 6 la_data_in[1]
port 157 nsew signal input
rlabel metal2 s 48042 0 48098 800 6 la_data_in[20]
port 158 nsew signal input
rlabel metal2 s 48870 0 48926 800 6 la_data_in[21]
port 159 nsew signal input
rlabel metal2 s 49790 0 49846 800 6 la_data_in[22]
port 160 nsew signal input
rlabel metal2 s 50618 0 50674 800 6 la_data_in[23]
port 161 nsew signal input
rlabel metal2 s 51538 0 51594 800 6 la_data_in[24]
port 162 nsew signal input
rlabel metal2 s 52366 0 52422 800 6 la_data_in[25]
port 163 nsew signal input
rlabel metal2 s 53286 0 53342 800 6 la_data_in[26]
port 164 nsew signal input
rlabel metal2 s 54114 0 54170 800 6 la_data_in[27]
port 165 nsew signal input
rlabel metal2 s 54942 0 54998 800 6 la_data_in[28]
port 166 nsew signal input
rlabel metal2 s 55862 0 55918 800 6 la_data_in[29]
port 167 nsew signal input
rlabel metal2 s 32402 0 32458 800 6 la_data_in[2]
port 168 nsew signal input
rlabel metal2 s 56690 0 56746 800 6 la_data_in[30]
port 169 nsew signal input
rlabel metal2 s 57610 0 57666 800 6 la_data_in[31]
port 170 nsew signal input
rlabel metal2 s 58438 0 58494 800 6 la_data_in[32]
port 171 nsew signal input
rlabel metal2 s 59358 0 59414 800 6 la_data_in[33]
port 172 nsew signal input
rlabel metal2 s 60186 0 60242 800 6 la_data_in[34]
port 173 nsew signal input
rlabel metal2 s 61014 0 61070 800 6 la_data_in[35]
port 174 nsew signal input
rlabel metal2 s 61934 0 61990 800 6 la_data_in[36]
port 175 nsew signal input
rlabel metal2 s 62762 0 62818 800 6 la_data_in[37]
port 176 nsew signal input
rlabel metal2 s 63682 0 63738 800 6 la_data_in[38]
port 177 nsew signal input
rlabel metal2 s 64510 0 64566 800 6 la_data_in[39]
port 178 nsew signal input
rlabel metal2 s 33322 0 33378 800 6 la_data_in[3]
port 179 nsew signal input
rlabel metal2 s 65430 0 65486 800 6 la_data_in[40]
port 180 nsew signal input
rlabel metal2 s 66258 0 66314 800 6 la_data_in[41]
port 181 nsew signal input
rlabel metal2 s 67086 0 67142 800 6 la_data_in[42]
port 182 nsew signal input
rlabel metal2 s 68006 0 68062 800 6 la_data_in[43]
port 183 nsew signal input
rlabel metal2 s 68834 0 68890 800 6 la_data_in[44]
port 184 nsew signal input
rlabel metal2 s 69754 0 69810 800 6 la_data_in[45]
port 185 nsew signal input
rlabel metal2 s 70582 0 70638 800 6 la_data_in[46]
port 186 nsew signal input
rlabel metal2 s 71502 0 71558 800 6 la_data_in[47]
port 187 nsew signal input
rlabel metal2 s 72330 0 72386 800 6 la_data_in[48]
port 188 nsew signal input
rlabel metal2 s 73158 0 73214 800 6 la_data_in[49]
port 189 nsew signal input
rlabel metal2 s 34150 0 34206 800 6 la_data_in[4]
port 190 nsew signal input
rlabel metal2 s 74078 0 74134 800 6 la_data_in[50]
port 191 nsew signal input
rlabel metal2 s 74906 0 74962 800 6 la_data_in[51]
port 192 nsew signal input
rlabel metal2 s 75826 0 75882 800 6 la_data_in[52]
port 193 nsew signal input
rlabel metal2 s 76654 0 76710 800 6 la_data_in[53]
port 194 nsew signal input
rlabel metal2 s 77574 0 77630 800 6 la_data_in[54]
port 195 nsew signal input
rlabel metal2 s 78402 0 78458 800 6 la_data_in[55]
port 196 nsew signal input
rlabel metal2 s 79230 0 79286 800 6 la_data_in[56]
port 197 nsew signal input
rlabel metal2 s 80150 0 80206 800 6 la_data_in[57]
port 198 nsew signal input
rlabel metal2 s 80978 0 81034 800 6 la_data_in[58]
port 199 nsew signal input
rlabel metal2 s 81898 0 81954 800 6 la_data_in[59]
port 200 nsew signal input
rlabel metal2 s 35070 0 35126 800 6 la_data_in[5]
port 201 nsew signal input
rlabel metal2 s 82726 0 82782 800 6 la_data_in[60]
port 202 nsew signal input
rlabel metal2 s 83646 0 83702 800 6 la_data_in[61]
port 203 nsew signal input
rlabel metal2 s 84474 0 84530 800 6 la_data_in[62]
port 204 nsew signal input
rlabel metal2 s 85302 0 85358 800 6 la_data_in[63]
port 205 nsew signal input
rlabel metal2 s 86222 0 86278 800 6 la_data_in[64]
port 206 nsew signal input
rlabel metal2 s 87050 0 87106 800 6 la_data_in[65]
port 207 nsew signal input
rlabel metal2 s 87970 0 88026 800 6 la_data_in[66]
port 208 nsew signal input
rlabel metal2 s 88798 0 88854 800 6 la_data_in[67]
port 209 nsew signal input
rlabel metal2 s 89718 0 89774 800 6 la_data_in[68]
port 210 nsew signal input
rlabel metal2 s 90546 0 90602 800 6 la_data_in[69]
port 211 nsew signal input
rlabel metal2 s 35898 0 35954 800 6 la_data_in[6]
port 212 nsew signal input
rlabel metal2 s 91374 0 91430 800 6 la_data_in[70]
port 213 nsew signal input
rlabel metal2 s 92294 0 92350 800 6 la_data_in[71]
port 214 nsew signal input
rlabel metal2 s 93122 0 93178 800 6 la_data_in[72]
port 215 nsew signal input
rlabel metal2 s 94042 0 94098 800 6 la_data_in[73]
port 216 nsew signal input
rlabel metal2 s 94870 0 94926 800 6 la_data_in[74]
port 217 nsew signal input
rlabel metal2 s 95698 0 95754 800 6 la_data_in[75]
port 218 nsew signal input
rlabel metal2 s 96618 0 96674 800 6 la_data_in[76]
port 219 nsew signal input
rlabel metal2 s 97446 0 97502 800 6 la_data_in[77]
port 220 nsew signal input
rlabel metal2 s 98366 0 98422 800 6 la_data_in[78]
port 221 nsew signal input
rlabel metal2 s 99194 0 99250 800 6 la_data_in[79]
port 222 nsew signal input
rlabel metal2 s 36818 0 36874 800 6 la_data_in[7]
port 223 nsew signal input
rlabel metal2 s 100114 0 100170 800 6 la_data_in[80]
port 224 nsew signal input
rlabel metal2 s 100942 0 100998 800 6 la_data_in[81]
port 225 nsew signal input
rlabel metal2 s 101770 0 101826 800 6 la_data_in[82]
port 226 nsew signal input
rlabel metal2 s 102690 0 102746 800 6 la_data_in[83]
port 227 nsew signal input
rlabel metal2 s 103518 0 103574 800 6 la_data_in[84]
port 228 nsew signal input
rlabel metal2 s 104438 0 104494 800 6 la_data_in[85]
port 229 nsew signal input
rlabel metal2 s 105266 0 105322 800 6 la_data_in[86]
port 230 nsew signal input
rlabel metal2 s 106186 0 106242 800 6 la_data_in[87]
port 231 nsew signal input
rlabel metal2 s 107014 0 107070 800 6 la_data_in[88]
port 232 nsew signal input
rlabel metal2 s 107842 0 107898 800 6 la_data_in[89]
port 233 nsew signal input
rlabel metal2 s 37646 0 37702 800 6 la_data_in[8]
port 234 nsew signal input
rlabel metal2 s 108762 0 108818 800 6 la_data_in[90]
port 235 nsew signal input
rlabel metal2 s 109590 0 109646 800 6 la_data_in[91]
port 236 nsew signal input
rlabel metal2 s 110510 0 110566 800 6 la_data_in[92]
port 237 nsew signal input
rlabel metal2 s 111338 0 111394 800 6 la_data_in[93]
port 238 nsew signal input
rlabel metal2 s 112258 0 112314 800 6 la_data_in[94]
port 239 nsew signal input
rlabel metal2 s 113086 0 113142 800 6 la_data_in[95]
port 240 nsew signal input
rlabel metal2 s 113914 0 113970 800 6 la_data_in[96]
port 241 nsew signal input
rlabel metal2 s 114834 0 114890 800 6 la_data_in[97]
port 242 nsew signal input
rlabel metal2 s 115662 0 115718 800 6 la_data_in[98]
port 243 nsew signal input
rlabel metal2 s 116582 0 116638 800 6 la_data_in[99]
port 244 nsew signal input
rlabel metal2 s 38474 0 38530 800 6 la_data_in[9]
port 245 nsew signal input
rlabel metal2 s 31022 0 31078 800 6 la_data_out[0]
port 246 nsew signal output
rlabel metal2 s 117686 0 117742 800 6 la_data_out[100]
port 247 nsew signal output
rlabel metal2 s 118606 0 118662 800 6 la_data_out[101]
port 248 nsew signal output
rlabel metal2 s 119434 0 119490 800 6 la_data_out[102]
port 249 nsew signal output
rlabel metal2 s 120354 0 120410 800 6 la_data_out[103]
port 250 nsew signal output
rlabel metal2 s 121182 0 121238 800 6 la_data_out[104]
port 251 nsew signal output
rlabel metal2 s 122010 0 122066 800 6 la_data_out[105]
port 252 nsew signal output
rlabel metal2 s 122930 0 122986 800 6 la_data_out[106]
port 253 nsew signal output
rlabel metal2 s 123758 0 123814 800 6 la_data_out[107]
port 254 nsew signal output
rlabel metal2 s 124678 0 124734 800 6 la_data_out[108]
port 255 nsew signal output
rlabel metal2 s 125506 0 125562 800 6 la_data_out[109]
port 256 nsew signal output
rlabel metal2 s 39670 0 39726 800 6 la_data_out[10]
port 257 nsew signal output
rlabel metal2 s 126426 0 126482 800 6 la_data_out[110]
port 258 nsew signal output
rlabel metal2 s 127254 0 127310 800 6 la_data_out[111]
port 259 nsew signal output
rlabel metal2 s 128082 0 128138 800 6 la_data_out[112]
port 260 nsew signal output
rlabel metal2 s 129002 0 129058 800 6 la_data_out[113]
port 261 nsew signal output
rlabel metal2 s 129830 0 129886 800 6 la_data_out[114]
port 262 nsew signal output
rlabel metal2 s 130750 0 130806 800 6 la_data_out[115]
port 263 nsew signal output
rlabel metal2 s 131578 0 131634 800 6 la_data_out[116]
port 264 nsew signal output
rlabel metal2 s 132498 0 132554 800 6 la_data_out[117]
port 265 nsew signal output
rlabel metal2 s 133326 0 133382 800 6 la_data_out[118]
port 266 nsew signal output
rlabel metal2 s 134154 0 134210 800 6 la_data_out[119]
port 267 nsew signal output
rlabel metal2 s 40498 0 40554 800 6 la_data_out[11]
port 268 nsew signal output
rlabel metal2 s 135074 0 135130 800 6 la_data_out[120]
port 269 nsew signal output
rlabel metal2 s 135902 0 135958 800 6 la_data_out[121]
port 270 nsew signal output
rlabel metal2 s 136822 0 136878 800 6 la_data_out[122]
port 271 nsew signal output
rlabel metal2 s 137650 0 137706 800 6 la_data_out[123]
port 272 nsew signal output
rlabel metal2 s 138570 0 138626 800 6 la_data_out[124]
port 273 nsew signal output
rlabel metal2 s 139398 0 139454 800 6 la_data_out[125]
port 274 nsew signal output
rlabel metal2 s 140226 0 140282 800 6 la_data_out[126]
port 275 nsew signal output
rlabel metal2 s 141146 0 141202 800 6 la_data_out[127]
port 276 nsew signal output
rlabel metal2 s 41418 0 41474 800 6 la_data_out[12]
port 277 nsew signal output
rlabel metal2 s 42246 0 42302 800 6 la_data_out[13]
port 278 nsew signal output
rlabel metal2 s 43166 0 43222 800 6 la_data_out[14]
port 279 nsew signal output
rlabel metal2 s 43994 0 44050 800 6 la_data_out[15]
port 280 nsew signal output
rlabel metal2 s 44914 0 44970 800 6 la_data_out[16]
port 281 nsew signal output
rlabel metal2 s 45742 0 45798 800 6 la_data_out[17]
port 282 nsew signal output
rlabel metal2 s 46570 0 46626 800 6 la_data_out[18]
port 283 nsew signal output
rlabel metal2 s 47490 0 47546 800 6 la_data_out[19]
port 284 nsew signal output
rlabel metal2 s 31850 0 31906 800 6 la_data_out[1]
port 285 nsew signal output
rlabel metal2 s 48318 0 48374 800 6 la_data_out[20]
port 286 nsew signal output
rlabel metal2 s 49238 0 49294 800 6 la_data_out[21]
port 287 nsew signal output
rlabel metal2 s 50066 0 50122 800 6 la_data_out[22]
port 288 nsew signal output
rlabel metal2 s 50894 0 50950 800 6 la_data_out[23]
port 289 nsew signal output
rlabel metal2 s 51814 0 51870 800 6 la_data_out[24]
port 290 nsew signal output
rlabel metal2 s 52642 0 52698 800 6 la_data_out[25]
port 291 nsew signal output
rlabel metal2 s 53562 0 53618 800 6 la_data_out[26]
port 292 nsew signal output
rlabel metal2 s 54390 0 54446 800 6 la_data_out[27]
port 293 nsew signal output
rlabel metal2 s 55310 0 55366 800 6 la_data_out[28]
port 294 nsew signal output
rlabel metal2 s 56138 0 56194 800 6 la_data_out[29]
port 295 nsew signal output
rlabel metal2 s 32770 0 32826 800 6 la_data_out[2]
port 296 nsew signal output
rlabel metal2 s 56966 0 57022 800 6 la_data_out[30]
port 297 nsew signal output
rlabel metal2 s 57886 0 57942 800 6 la_data_out[31]
port 298 nsew signal output
rlabel metal2 s 58714 0 58770 800 6 la_data_out[32]
port 299 nsew signal output
rlabel metal2 s 59634 0 59690 800 6 la_data_out[33]
port 300 nsew signal output
rlabel metal2 s 60462 0 60518 800 6 la_data_out[34]
port 301 nsew signal output
rlabel metal2 s 61382 0 61438 800 6 la_data_out[35]
port 302 nsew signal output
rlabel metal2 s 62210 0 62266 800 6 la_data_out[36]
port 303 nsew signal output
rlabel metal2 s 63038 0 63094 800 6 la_data_out[37]
port 304 nsew signal output
rlabel metal2 s 63958 0 64014 800 6 la_data_out[38]
port 305 nsew signal output
rlabel metal2 s 64786 0 64842 800 6 la_data_out[39]
port 306 nsew signal output
rlabel metal2 s 33598 0 33654 800 6 la_data_out[3]
port 307 nsew signal output
rlabel metal2 s 65706 0 65762 800 6 la_data_out[40]
port 308 nsew signal output
rlabel metal2 s 66534 0 66590 800 6 la_data_out[41]
port 309 nsew signal output
rlabel metal2 s 67454 0 67510 800 6 la_data_out[42]
port 310 nsew signal output
rlabel metal2 s 68282 0 68338 800 6 la_data_out[43]
port 311 nsew signal output
rlabel metal2 s 69110 0 69166 800 6 la_data_out[44]
port 312 nsew signal output
rlabel metal2 s 70030 0 70086 800 6 la_data_out[45]
port 313 nsew signal output
rlabel metal2 s 70858 0 70914 800 6 la_data_out[46]
port 314 nsew signal output
rlabel metal2 s 71778 0 71834 800 6 la_data_out[47]
port 315 nsew signal output
rlabel metal2 s 72606 0 72662 800 6 la_data_out[48]
port 316 nsew signal output
rlabel metal2 s 73526 0 73582 800 6 la_data_out[49]
port 317 nsew signal output
rlabel metal2 s 34426 0 34482 800 6 la_data_out[4]
port 318 nsew signal output
rlabel metal2 s 74354 0 74410 800 6 la_data_out[50]
port 319 nsew signal output
rlabel metal2 s 75182 0 75238 800 6 la_data_out[51]
port 320 nsew signal output
rlabel metal2 s 76102 0 76158 800 6 la_data_out[52]
port 321 nsew signal output
rlabel metal2 s 76930 0 76986 800 6 la_data_out[53]
port 322 nsew signal output
rlabel metal2 s 77850 0 77906 800 6 la_data_out[54]
port 323 nsew signal output
rlabel metal2 s 78678 0 78734 800 6 la_data_out[55]
port 324 nsew signal output
rlabel metal2 s 79598 0 79654 800 6 la_data_out[56]
port 325 nsew signal output
rlabel metal2 s 80426 0 80482 800 6 la_data_out[57]
port 326 nsew signal output
rlabel metal2 s 81254 0 81310 800 6 la_data_out[58]
port 327 nsew signal output
rlabel metal2 s 82174 0 82230 800 6 la_data_out[59]
port 328 nsew signal output
rlabel metal2 s 35346 0 35402 800 6 la_data_out[5]
port 329 nsew signal output
rlabel metal2 s 83002 0 83058 800 6 la_data_out[60]
port 330 nsew signal output
rlabel metal2 s 83922 0 83978 800 6 la_data_out[61]
port 331 nsew signal output
rlabel metal2 s 84750 0 84806 800 6 la_data_out[62]
port 332 nsew signal output
rlabel metal2 s 85670 0 85726 800 6 la_data_out[63]
port 333 nsew signal output
rlabel metal2 s 86498 0 86554 800 6 la_data_out[64]
port 334 nsew signal output
rlabel metal2 s 87326 0 87382 800 6 la_data_out[65]
port 335 nsew signal output
rlabel metal2 s 88246 0 88302 800 6 la_data_out[66]
port 336 nsew signal output
rlabel metal2 s 89074 0 89130 800 6 la_data_out[67]
port 337 nsew signal output
rlabel metal2 s 89994 0 90050 800 6 la_data_out[68]
port 338 nsew signal output
rlabel metal2 s 90822 0 90878 800 6 la_data_out[69]
port 339 nsew signal output
rlabel metal2 s 36174 0 36230 800 6 la_data_out[6]
port 340 nsew signal output
rlabel metal2 s 91742 0 91798 800 6 la_data_out[70]
port 341 nsew signal output
rlabel metal2 s 92570 0 92626 800 6 la_data_out[71]
port 342 nsew signal output
rlabel metal2 s 93398 0 93454 800 6 la_data_out[72]
port 343 nsew signal output
rlabel metal2 s 94318 0 94374 800 6 la_data_out[73]
port 344 nsew signal output
rlabel metal2 s 95146 0 95202 800 6 la_data_out[74]
port 345 nsew signal output
rlabel metal2 s 96066 0 96122 800 6 la_data_out[75]
port 346 nsew signal output
rlabel metal2 s 96894 0 96950 800 6 la_data_out[76]
port 347 nsew signal output
rlabel metal2 s 97722 0 97778 800 6 la_data_out[77]
port 348 nsew signal output
rlabel metal2 s 98642 0 98698 800 6 la_data_out[78]
port 349 nsew signal output
rlabel metal2 s 99470 0 99526 800 6 la_data_out[79]
port 350 nsew signal output
rlabel metal2 s 37094 0 37150 800 6 la_data_out[7]
port 351 nsew signal output
rlabel metal2 s 100390 0 100446 800 6 la_data_out[80]
port 352 nsew signal output
rlabel metal2 s 101218 0 101274 800 6 la_data_out[81]
port 353 nsew signal output
rlabel metal2 s 102138 0 102194 800 6 la_data_out[82]
port 354 nsew signal output
rlabel metal2 s 102966 0 103022 800 6 la_data_out[83]
port 355 nsew signal output
rlabel metal2 s 103794 0 103850 800 6 la_data_out[84]
port 356 nsew signal output
rlabel metal2 s 104714 0 104770 800 6 la_data_out[85]
port 357 nsew signal output
rlabel metal2 s 105542 0 105598 800 6 la_data_out[86]
port 358 nsew signal output
rlabel metal2 s 106462 0 106518 800 6 la_data_out[87]
port 359 nsew signal output
rlabel metal2 s 107290 0 107346 800 6 la_data_out[88]
port 360 nsew signal output
rlabel metal2 s 108210 0 108266 800 6 la_data_out[89]
port 361 nsew signal output
rlabel metal2 s 37922 0 37978 800 6 la_data_out[8]
port 362 nsew signal output
rlabel metal2 s 109038 0 109094 800 6 la_data_out[90]
port 363 nsew signal output
rlabel metal2 s 109866 0 109922 800 6 la_data_out[91]
port 364 nsew signal output
rlabel metal2 s 110786 0 110842 800 6 la_data_out[92]
port 365 nsew signal output
rlabel metal2 s 111614 0 111670 800 6 la_data_out[93]
port 366 nsew signal output
rlabel metal2 s 112534 0 112590 800 6 la_data_out[94]
port 367 nsew signal output
rlabel metal2 s 113362 0 113418 800 6 la_data_out[95]
port 368 nsew signal output
rlabel metal2 s 114282 0 114338 800 6 la_data_out[96]
port 369 nsew signal output
rlabel metal2 s 115110 0 115166 800 6 la_data_out[97]
port 370 nsew signal output
rlabel metal2 s 115938 0 115994 800 6 la_data_out[98]
port 371 nsew signal output
rlabel metal2 s 116858 0 116914 800 6 la_data_out[99]
port 372 nsew signal output
rlabel metal2 s 38842 0 38898 800 6 la_data_out[9]
port 373 nsew signal output
rlabel metal2 s 31298 0 31354 800 6 la_oenb[0]
port 374 nsew signal input
rlabel metal2 s 117962 0 118018 800 6 la_oenb[100]
port 375 nsew signal input
rlabel metal2 s 118882 0 118938 800 6 la_oenb[101]
port 376 nsew signal input
rlabel metal2 s 119710 0 119766 800 6 la_oenb[102]
port 377 nsew signal input
rlabel metal2 s 120630 0 120686 800 6 la_oenb[103]
port 378 nsew signal input
rlabel metal2 s 121458 0 121514 800 6 la_oenb[104]
port 379 nsew signal input
rlabel metal2 s 122378 0 122434 800 6 la_oenb[105]
port 380 nsew signal input
rlabel metal2 s 123206 0 123262 800 6 la_oenb[106]
port 381 nsew signal input
rlabel metal2 s 124034 0 124090 800 6 la_oenb[107]
port 382 nsew signal input
rlabel metal2 s 124954 0 125010 800 6 la_oenb[108]
port 383 nsew signal input
rlabel metal2 s 125782 0 125838 800 6 la_oenb[109]
port 384 nsew signal input
rlabel metal2 s 39946 0 40002 800 6 la_oenb[10]
port 385 nsew signal input
rlabel metal2 s 126702 0 126758 800 6 la_oenb[110]
port 386 nsew signal input
rlabel metal2 s 127530 0 127586 800 6 la_oenb[111]
port 387 nsew signal input
rlabel metal2 s 128450 0 128506 800 6 la_oenb[112]
port 388 nsew signal input
rlabel metal2 s 129278 0 129334 800 6 la_oenb[113]
port 389 nsew signal input
rlabel metal2 s 130106 0 130162 800 6 la_oenb[114]
port 390 nsew signal input
rlabel metal2 s 131026 0 131082 800 6 la_oenb[115]
port 391 nsew signal input
rlabel metal2 s 131854 0 131910 800 6 la_oenb[116]
port 392 nsew signal input
rlabel metal2 s 132774 0 132830 800 6 la_oenb[117]
port 393 nsew signal input
rlabel metal2 s 133602 0 133658 800 6 la_oenb[118]
port 394 nsew signal input
rlabel metal2 s 134522 0 134578 800 6 la_oenb[119]
port 395 nsew signal input
rlabel metal2 s 40866 0 40922 800 6 la_oenb[11]
port 396 nsew signal input
rlabel metal2 s 135350 0 135406 800 6 la_oenb[120]
port 397 nsew signal input
rlabel metal2 s 136178 0 136234 800 6 la_oenb[121]
port 398 nsew signal input
rlabel metal2 s 137098 0 137154 800 6 la_oenb[122]
port 399 nsew signal input
rlabel metal2 s 137926 0 137982 800 6 la_oenb[123]
port 400 nsew signal input
rlabel metal2 s 138846 0 138902 800 6 la_oenb[124]
port 401 nsew signal input
rlabel metal2 s 139674 0 139730 800 6 la_oenb[125]
port 402 nsew signal input
rlabel metal2 s 140594 0 140650 800 6 la_oenb[126]
port 403 nsew signal input
rlabel metal2 s 141422 0 141478 800 6 la_oenb[127]
port 404 nsew signal input
rlabel metal2 s 41694 0 41750 800 6 la_oenb[12]
port 405 nsew signal input
rlabel metal2 s 42522 0 42578 800 6 la_oenb[13]
port 406 nsew signal input
rlabel metal2 s 43442 0 43498 800 6 la_oenb[14]
port 407 nsew signal input
rlabel metal2 s 44270 0 44326 800 6 la_oenb[15]
port 408 nsew signal input
rlabel metal2 s 45190 0 45246 800 6 la_oenb[16]
port 409 nsew signal input
rlabel metal2 s 46018 0 46074 800 6 la_oenb[17]
port 410 nsew signal input
rlabel metal2 s 46938 0 46994 800 6 la_oenb[18]
port 411 nsew signal input
rlabel metal2 s 47766 0 47822 800 6 la_oenb[19]
port 412 nsew signal input
rlabel metal2 s 32126 0 32182 800 6 la_oenb[1]
port 413 nsew signal input
rlabel metal2 s 48594 0 48650 800 6 la_oenb[20]
port 414 nsew signal input
rlabel metal2 s 49514 0 49570 800 6 la_oenb[21]
port 415 nsew signal input
rlabel metal2 s 50342 0 50398 800 6 la_oenb[22]
port 416 nsew signal input
rlabel metal2 s 51262 0 51318 800 6 la_oenb[23]
port 417 nsew signal input
rlabel metal2 s 52090 0 52146 800 6 la_oenb[24]
port 418 nsew signal input
rlabel metal2 s 52918 0 52974 800 6 la_oenb[25]
port 419 nsew signal input
rlabel metal2 s 53838 0 53894 800 6 la_oenb[26]
port 420 nsew signal input
rlabel metal2 s 54666 0 54722 800 6 la_oenb[27]
port 421 nsew signal input
rlabel metal2 s 55586 0 55642 800 6 la_oenb[28]
port 422 nsew signal input
rlabel metal2 s 56414 0 56470 800 6 la_oenb[29]
port 423 nsew signal input
rlabel metal2 s 33046 0 33102 800 6 la_oenb[2]
port 424 nsew signal input
rlabel metal2 s 57334 0 57390 800 6 la_oenb[30]
port 425 nsew signal input
rlabel metal2 s 58162 0 58218 800 6 la_oenb[31]
port 426 nsew signal input
rlabel metal2 s 58990 0 59046 800 6 la_oenb[32]
port 427 nsew signal input
rlabel metal2 s 59910 0 59966 800 6 la_oenb[33]
port 428 nsew signal input
rlabel metal2 s 60738 0 60794 800 6 la_oenb[34]
port 429 nsew signal input
rlabel metal2 s 61658 0 61714 800 6 la_oenb[35]
port 430 nsew signal input
rlabel metal2 s 62486 0 62542 800 6 la_oenb[36]
port 431 nsew signal input
rlabel metal2 s 63406 0 63462 800 6 la_oenb[37]
port 432 nsew signal input
rlabel metal2 s 64234 0 64290 800 6 la_oenb[38]
port 433 nsew signal input
rlabel metal2 s 65062 0 65118 800 6 la_oenb[39]
port 434 nsew signal input
rlabel metal2 s 33874 0 33930 800 6 la_oenb[3]
port 435 nsew signal input
rlabel metal2 s 65982 0 66038 800 6 la_oenb[40]
port 436 nsew signal input
rlabel metal2 s 66810 0 66866 800 6 la_oenb[41]
port 437 nsew signal input
rlabel metal2 s 67730 0 67786 800 6 la_oenb[42]
port 438 nsew signal input
rlabel metal2 s 68558 0 68614 800 6 la_oenb[43]
port 439 nsew signal input
rlabel metal2 s 69478 0 69534 800 6 la_oenb[44]
port 440 nsew signal input
rlabel metal2 s 70306 0 70362 800 6 la_oenb[45]
port 441 nsew signal input
rlabel metal2 s 71134 0 71190 800 6 la_oenb[46]
port 442 nsew signal input
rlabel metal2 s 72054 0 72110 800 6 la_oenb[47]
port 443 nsew signal input
rlabel metal2 s 72882 0 72938 800 6 la_oenb[48]
port 444 nsew signal input
rlabel metal2 s 73802 0 73858 800 6 la_oenb[49]
port 445 nsew signal input
rlabel metal2 s 34794 0 34850 800 6 la_oenb[4]
port 446 nsew signal input
rlabel metal2 s 74630 0 74686 800 6 la_oenb[50]
port 447 nsew signal input
rlabel metal2 s 75550 0 75606 800 6 la_oenb[51]
port 448 nsew signal input
rlabel metal2 s 76378 0 76434 800 6 la_oenb[52]
port 449 nsew signal input
rlabel metal2 s 77206 0 77262 800 6 la_oenb[53]
port 450 nsew signal input
rlabel metal2 s 78126 0 78182 800 6 la_oenb[54]
port 451 nsew signal input
rlabel metal2 s 78954 0 79010 800 6 la_oenb[55]
port 452 nsew signal input
rlabel metal2 s 79874 0 79930 800 6 la_oenb[56]
port 453 nsew signal input
rlabel metal2 s 80702 0 80758 800 6 la_oenb[57]
port 454 nsew signal input
rlabel metal2 s 81622 0 81678 800 6 la_oenb[58]
port 455 nsew signal input
rlabel metal2 s 82450 0 82506 800 6 la_oenb[59]
port 456 nsew signal input
rlabel metal2 s 35622 0 35678 800 6 la_oenb[5]
port 457 nsew signal input
rlabel metal2 s 83278 0 83334 800 6 la_oenb[60]
port 458 nsew signal input
rlabel metal2 s 84198 0 84254 800 6 la_oenb[61]
port 459 nsew signal input
rlabel metal2 s 85026 0 85082 800 6 la_oenb[62]
port 460 nsew signal input
rlabel metal2 s 85946 0 86002 800 6 la_oenb[63]
port 461 nsew signal input
rlabel metal2 s 86774 0 86830 800 6 la_oenb[64]
port 462 nsew signal input
rlabel metal2 s 87694 0 87750 800 6 la_oenb[65]
port 463 nsew signal input
rlabel metal2 s 88522 0 88578 800 6 la_oenb[66]
port 464 nsew signal input
rlabel metal2 s 89350 0 89406 800 6 la_oenb[67]
port 465 nsew signal input
rlabel metal2 s 90270 0 90326 800 6 la_oenb[68]
port 466 nsew signal input
rlabel metal2 s 91098 0 91154 800 6 la_oenb[69]
port 467 nsew signal input
rlabel metal2 s 36450 0 36506 800 6 la_oenb[6]
port 468 nsew signal input
rlabel metal2 s 92018 0 92074 800 6 la_oenb[70]
port 469 nsew signal input
rlabel metal2 s 92846 0 92902 800 6 la_oenb[71]
port 470 nsew signal input
rlabel metal2 s 93766 0 93822 800 6 la_oenb[72]
port 471 nsew signal input
rlabel metal2 s 94594 0 94650 800 6 la_oenb[73]
port 472 nsew signal input
rlabel metal2 s 95422 0 95478 800 6 la_oenb[74]
port 473 nsew signal input
rlabel metal2 s 96342 0 96398 800 6 la_oenb[75]
port 474 nsew signal input
rlabel metal2 s 97170 0 97226 800 6 la_oenb[76]
port 475 nsew signal input
rlabel metal2 s 98090 0 98146 800 6 la_oenb[77]
port 476 nsew signal input
rlabel metal2 s 98918 0 98974 800 6 la_oenb[78]
port 477 nsew signal input
rlabel metal2 s 99746 0 99802 800 6 la_oenb[79]
port 478 nsew signal input
rlabel metal2 s 37370 0 37426 800 6 la_oenb[7]
port 479 nsew signal input
rlabel metal2 s 100666 0 100722 800 6 la_oenb[80]
port 480 nsew signal input
rlabel metal2 s 101494 0 101550 800 6 la_oenb[81]
port 481 nsew signal input
rlabel metal2 s 102414 0 102470 800 6 la_oenb[82]
port 482 nsew signal input
rlabel metal2 s 103242 0 103298 800 6 la_oenb[83]
port 483 nsew signal input
rlabel metal2 s 104162 0 104218 800 6 la_oenb[84]
port 484 nsew signal input
rlabel metal2 s 104990 0 105046 800 6 la_oenb[85]
port 485 nsew signal input
rlabel metal2 s 105818 0 105874 800 6 la_oenb[86]
port 486 nsew signal input
rlabel metal2 s 106738 0 106794 800 6 la_oenb[87]
port 487 nsew signal input
rlabel metal2 s 107566 0 107622 800 6 la_oenb[88]
port 488 nsew signal input
rlabel metal2 s 108486 0 108542 800 6 la_oenb[89]
port 489 nsew signal input
rlabel metal2 s 38198 0 38254 800 6 la_oenb[8]
port 490 nsew signal input
rlabel metal2 s 109314 0 109370 800 6 la_oenb[90]
port 491 nsew signal input
rlabel metal2 s 110234 0 110290 800 6 la_oenb[91]
port 492 nsew signal input
rlabel metal2 s 111062 0 111118 800 6 la_oenb[92]
port 493 nsew signal input
rlabel metal2 s 111890 0 111946 800 6 la_oenb[93]
port 494 nsew signal input
rlabel metal2 s 112810 0 112866 800 6 la_oenb[94]
port 495 nsew signal input
rlabel metal2 s 113638 0 113694 800 6 la_oenb[95]
port 496 nsew signal input
rlabel metal2 s 114558 0 114614 800 6 la_oenb[96]
port 497 nsew signal input
rlabel metal2 s 115386 0 115442 800 6 la_oenb[97]
port 498 nsew signal input
rlabel metal2 s 116306 0 116362 800 6 la_oenb[98]
port 499 nsew signal input
rlabel metal2 s 117134 0 117190 800 6 la_oenb[99]
port 500 nsew signal input
rlabel metal2 s 39118 0 39174 800 6 la_oenb[9]
port 501 nsew signal input
rlabel metal4 s 4208 2128 4528 142032 6 vccd1
port 502 nsew power input
rlabel metal4 s 34928 2128 35248 142032 6 vccd1
port 502 nsew power input
rlabel metal4 s 65648 2128 65968 142032 6 vccd1
port 502 nsew power input
rlabel metal4 s 96368 2128 96688 142032 6 vccd1
port 502 nsew power input
rlabel metal4 s 127088 2128 127408 142032 6 vccd1
port 502 nsew power input
rlabel metal4 s 19568 2128 19888 142032 6 vssd1
port 503 nsew ground input
rlabel metal4 s 50288 2128 50608 142032 6 vssd1
port 503 nsew ground input
rlabel metal4 s 81008 2128 81328 142032 6 vssd1
port 503 nsew ground input
rlabel metal4 s 111728 2128 112048 142032 6 vssd1
port 503 nsew ground input
rlabel metal2 s 110 0 166 800 6 wb_clk_i
port 504 nsew signal input
rlabel metal2 s 386 0 442 800 6 wb_rst_i
port 505 nsew signal input
rlabel metal2 s 662 0 718 800 6 wbs_ack_o
port 506 nsew signal output
rlabel metal2 s 1766 0 1822 800 6 wbs_adr_i[0]
port 507 nsew signal input
rlabel metal2 s 11610 0 11666 800 6 wbs_adr_i[10]
port 508 nsew signal input
rlabel metal2 s 12530 0 12586 800 6 wbs_adr_i[11]
port 509 nsew signal input
rlabel metal2 s 13358 0 13414 800 6 wbs_adr_i[12]
port 510 nsew signal input
rlabel metal2 s 14186 0 14242 800 6 wbs_adr_i[13]
port 511 nsew signal input
rlabel metal2 s 15106 0 15162 800 6 wbs_adr_i[14]
port 512 nsew signal input
rlabel metal2 s 15934 0 15990 800 6 wbs_adr_i[15]
port 513 nsew signal input
rlabel metal2 s 16854 0 16910 800 6 wbs_adr_i[16]
port 514 nsew signal input
rlabel metal2 s 17682 0 17738 800 6 wbs_adr_i[17]
port 515 nsew signal input
rlabel metal2 s 18602 0 18658 800 6 wbs_adr_i[18]
port 516 nsew signal input
rlabel metal2 s 19430 0 19486 800 6 wbs_adr_i[19]
port 517 nsew signal input
rlabel metal2 s 2962 0 3018 800 6 wbs_adr_i[1]
port 518 nsew signal input
rlabel metal2 s 20258 0 20314 800 6 wbs_adr_i[20]
port 519 nsew signal input
rlabel metal2 s 21178 0 21234 800 6 wbs_adr_i[21]
port 520 nsew signal input
rlabel metal2 s 22006 0 22062 800 6 wbs_adr_i[22]
port 521 nsew signal input
rlabel metal2 s 22926 0 22982 800 6 wbs_adr_i[23]
port 522 nsew signal input
rlabel metal2 s 23754 0 23810 800 6 wbs_adr_i[24]
port 523 nsew signal input
rlabel metal2 s 24674 0 24730 800 6 wbs_adr_i[25]
port 524 nsew signal input
rlabel metal2 s 25502 0 25558 800 6 wbs_adr_i[26]
port 525 nsew signal input
rlabel metal2 s 26330 0 26386 800 6 wbs_adr_i[27]
port 526 nsew signal input
rlabel metal2 s 27250 0 27306 800 6 wbs_adr_i[28]
port 527 nsew signal input
rlabel metal2 s 28078 0 28134 800 6 wbs_adr_i[29]
port 528 nsew signal input
rlabel metal2 s 4066 0 4122 800 6 wbs_adr_i[2]
port 529 nsew signal input
rlabel metal2 s 28998 0 29054 800 6 wbs_adr_i[30]
port 530 nsew signal input
rlabel metal2 s 29826 0 29882 800 6 wbs_adr_i[31]
port 531 nsew signal input
rlabel metal2 s 5262 0 5318 800 6 wbs_adr_i[3]
port 532 nsew signal input
rlabel metal2 s 6458 0 6514 800 6 wbs_adr_i[4]
port 533 nsew signal input
rlabel metal2 s 7286 0 7342 800 6 wbs_adr_i[5]
port 534 nsew signal input
rlabel metal2 s 8114 0 8170 800 6 wbs_adr_i[6]
port 535 nsew signal input
rlabel metal2 s 9034 0 9090 800 6 wbs_adr_i[7]
port 536 nsew signal input
rlabel metal2 s 9862 0 9918 800 6 wbs_adr_i[8]
port 537 nsew signal input
rlabel metal2 s 10782 0 10838 800 6 wbs_adr_i[9]
port 538 nsew signal input
rlabel metal2 s 938 0 994 800 6 wbs_cyc_i
port 539 nsew signal input
rlabel metal2 s 2042 0 2098 800 6 wbs_dat_i[0]
port 540 nsew signal input
rlabel metal2 s 11886 0 11942 800 6 wbs_dat_i[10]
port 541 nsew signal input
rlabel metal2 s 12806 0 12862 800 6 wbs_dat_i[11]
port 542 nsew signal input
rlabel metal2 s 13634 0 13690 800 6 wbs_dat_i[12]
port 543 nsew signal input
rlabel metal2 s 14554 0 14610 800 6 wbs_dat_i[13]
port 544 nsew signal input
rlabel metal2 s 15382 0 15438 800 6 wbs_dat_i[14]
port 545 nsew signal input
rlabel metal2 s 16210 0 16266 800 6 wbs_dat_i[15]
port 546 nsew signal input
rlabel metal2 s 17130 0 17186 800 6 wbs_dat_i[16]
port 547 nsew signal input
rlabel metal2 s 17958 0 18014 800 6 wbs_dat_i[17]
port 548 nsew signal input
rlabel metal2 s 18878 0 18934 800 6 wbs_dat_i[18]
port 549 nsew signal input
rlabel metal2 s 19706 0 19762 800 6 wbs_dat_i[19]
port 550 nsew signal input
rlabel metal2 s 3238 0 3294 800 6 wbs_dat_i[1]
port 551 nsew signal input
rlabel metal2 s 20626 0 20682 800 6 wbs_dat_i[20]
port 552 nsew signal input
rlabel metal2 s 21454 0 21510 800 6 wbs_dat_i[21]
port 553 nsew signal input
rlabel metal2 s 22282 0 22338 800 6 wbs_dat_i[22]
port 554 nsew signal input
rlabel metal2 s 23202 0 23258 800 6 wbs_dat_i[23]
port 555 nsew signal input
rlabel metal2 s 24030 0 24086 800 6 wbs_dat_i[24]
port 556 nsew signal input
rlabel metal2 s 24950 0 25006 800 6 wbs_dat_i[25]
port 557 nsew signal input
rlabel metal2 s 25778 0 25834 800 6 wbs_dat_i[26]
port 558 nsew signal input
rlabel metal2 s 26698 0 26754 800 6 wbs_dat_i[27]
port 559 nsew signal input
rlabel metal2 s 27526 0 27582 800 6 wbs_dat_i[28]
port 560 nsew signal input
rlabel metal2 s 28354 0 28410 800 6 wbs_dat_i[29]
port 561 nsew signal input
rlabel metal2 s 4434 0 4490 800 6 wbs_dat_i[2]
port 562 nsew signal input
rlabel metal2 s 29274 0 29330 800 6 wbs_dat_i[30]
port 563 nsew signal input
rlabel metal2 s 30102 0 30158 800 6 wbs_dat_i[31]
port 564 nsew signal input
rlabel metal2 s 5538 0 5594 800 6 wbs_dat_i[3]
port 565 nsew signal input
rlabel metal2 s 6734 0 6790 800 6 wbs_dat_i[4]
port 566 nsew signal input
rlabel metal2 s 7562 0 7618 800 6 wbs_dat_i[5]
port 567 nsew signal input
rlabel metal2 s 8482 0 8538 800 6 wbs_dat_i[6]
port 568 nsew signal input
rlabel metal2 s 9310 0 9366 800 6 wbs_dat_i[7]
port 569 nsew signal input
rlabel metal2 s 10138 0 10194 800 6 wbs_dat_i[8]
port 570 nsew signal input
rlabel metal2 s 11058 0 11114 800 6 wbs_dat_i[9]
port 571 nsew signal input
rlabel metal2 s 2410 0 2466 800 6 wbs_dat_o[0]
port 572 nsew signal output
rlabel metal2 s 12162 0 12218 800 6 wbs_dat_o[10]
port 573 nsew signal output
rlabel metal2 s 13082 0 13138 800 6 wbs_dat_o[11]
port 574 nsew signal output
rlabel metal2 s 13910 0 13966 800 6 wbs_dat_o[12]
port 575 nsew signal output
rlabel metal2 s 14830 0 14886 800 6 wbs_dat_o[13]
port 576 nsew signal output
rlabel metal2 s 15658 0 15714 800 6 wbs_dat_o[14]
port 577 nsew signal output
rlabel metal2 s 16578 0 16634 800 6 wbs_dat_o[15]
port 578 nsew signal output
rlabel metal2 s 17406 0 17462 800 6 wbs_dat_o[16]
port 579 nsew signal output
rlabel metal2 s 18234 0 18290 800 6 wbs_dat_o[17]
port 580 nsew signal output
rlabel metal2 s 19154 0 19210 800 6 wbs_dat_o[18]
port 581 nsew signal output
rlabel metal2 s 19982 0 20038 800 6 wbs_dat_o[19]
port 582 nsew signal output
rlabel metal2 s 3514 0 3570 800 6 wbs_dat_o[1]
port 583 nsew signal output
rlabel metal2 s 20902 0 20958 800 6 wbs_dat_o[20]
port 584 nsew signal output
rlabel metal2 s 21730 0 21786 800 6 wbs_dat_o[21]
port 585 nsew signal output
rlabel metal2 s 22650 0 22706 800 6 wbs_dat_o[22]
port 586 nsew signal output
rlabel metal2 s 23478 0 23534 800 6 wbs_dat_o[23]
port 587 nsew signal output
rlabel metal2 s 24306 0 24362 800 6 wbs_dat_o[24]
port 588 nsew signal output
rlabel metal2 s 25226 0 25282 800 6 wbs_dat_o[25]
port 589 nsew signal output
rlabel metal2 s 26054 0 26110 800 6 wbs_dat_o[26]
port 590 nsew signal output
rlabel metal2 s 26974 0 27030 800 6 wbs_dat_o[27]
port 591 nsew signal output
rlabel metal2 s 27802 0 27858 800 6 wbs_dat_o[28]
port 592 nsew signal output
rlabel metal2 s 28722 0 28778 800 6 wbs_dat_o[29]
port 593 nsew signal output
rlabel metal2 s 4710 0 4766 800 6 wbs_dat_o[2]
port 594 nsew signal output
rlabel metal2 s 29550 0 29606 800 6 wbs_dat_o[30]
port 595 nsew signal output
rlabel metal2 s 30378 0 30434 800 6 wbs_dat_o[31]
port 596 nsew signal output
rlabel metal2 s 5814 0 5870 800 6 wbs_dat_o[3]
port 597 nsew signal output
rlabel metal2 s 7010 0 7066 800 6 wbs_dat_o[4]
port 598 nsew signal output
rlabel metal2 s 7838 0 7894 800 6 wbs_dat_o[5]
port 599 nsew signal output
rlabel metal2 s 8758 0 8814 800 6 wbs_dat_o[6]
port 600 nsew signal output
rlabel metal2 s 9586 0 9642 800 6 wbs_dat_o[7]
port 601 nsew signal output
rlabel metal2 s 10506 0 10562 800 6 wbs_dat_o[8]
port 602 nsew signal output
rlabel metal2 s 11334 0 11390 800 6 wbs_dat_o[9]
port 603 nsew signal output
rlabel metal2 s 2686 0 2742 800 6 wbs_sel_i[0]
port 604 nsew signal input
rlabel metal2 s 3790 0 3846 800 6 wbs_sel_i[1]
port 605 nsew signal input
rlabel metal2 s 4986 0 5042 800 6 wbs_sel_i[2]
port 606 nsew signal input
rlabel metal2 s 6090 0 6146 800 6 wbs_sel_i[3]
port 607 nsew signal input
rlabel metal2 s 1214 0 1270 800 6 wbs_stb_i
port 608 nsew signal input
rlabel metal2 s 1490 0 1546 800 6 wbs_we_i
port 609 nsew signal input
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 142476 144620
string LEFview TRUE
string GDS_FILE /project/openlane/user_proj_example/runs/user_proj_example/results/magic/user_proj_example.gds
string GDS_END 59836198
string GDS_START 875772
<< end >>

