module sbox4(
    input [5:0] i_data,
    output reg [3:0] o_data
);



    always@(i_data) begin
        case(i_data)
            6'b000000: o_data = 4'b0111; // (0, 0) = 7
            6'b000001: o_data = 4'b1101; // (0, 1) = 13
            6'b000010: o_data = 4'b1101; // (1, 0) = 13
            6'b000011: o_data = 4'b1000; // (1, 1) = 8
            6'b000100: o_data = 4'b1110; // (2, 0) = 14
            6'b000101: o_data = 4'b1011; // (2, 1) = 11
            6'b000110: o_data = 4'b0011; // (3, 0) = 3
            6'b000111: o_data = 4'b0101; // (3, 1) = 5
            6'b001000: o_data = 4'b0000; // (4, 0) = 0
            6'b001001: o_data = 4'b0110; // (4, 1) = 6
            6'b001010: o_data = 4'b0110; // (5, 0) = 6
            6'b001011: o_data = 4'b1111; // (5, 1) = 15
            6'b001100: o_data = 4'b1001; // (6, 0) = 9
            6'b001101: o_data = 4'b0000; // (6, 1) = 0
            6'b001110: o_data = 4'b1010; // (7, 0) = 10
            6'b001111: o_data = 4'b0011; // (7, 1) = 3
            6'b010000: o_data = 4'b0001; // (8, 0) = 1
            6'b010001: o_data = 4'b0100; // (8, 1) = 4
            6'b010010: o_data = 4'b0010; // (9, 0) = 2
            6'b010011: o_data = 4'b0111; // (9, 1) = 7
            6'b010100: o_data = 4'b1000; // (10, 0) = 8
            6'b010101: o_data = 4'b0010; // (10, 1) = 2
            6'b010110: o_data = 4'b0101; // (11, 0) = 5
            6'b010111: o_data = 4'b1100; // (11, 1) = 12
            6'b011000: o_data = 4'b1011; // (12, 0) = 11
            6'b011001: o_data = 4'b0001; // (12, 1) = 1
            6'b011010: o_data = 4'b1100; // (13, 0) = 12
            6'b011011: o_data = 4'b1010; // (13, 1) = 10
            6'b011100: o_data = 4'b0100; // (14, 0) = 4
            6'b011101: o_data = 4'b1110; // (14, 1) = 14
            6'b011110: o_data = 4'b1111; // (15, 0) = 15
            6'b011111: o_data = 4'b1001; // (15, 1) = 9
            6'b100000: o_data = 4'b1010; // (0, 2) = 10
            6'b100001: o_data = 4'b0011; // (0, 3) = 3
            6'b100010: o_data = 4'b0110; // (1, 2) = 6
            6'b100011: o_data = 4'b1111; // (1, 3) = 15
            6'b100100: o_data = 4'b1001; // (2, 2) = 9
            6'b100101: o_data = 4'b0000; // (2, 3) = 0
            6'b100110: o_data = 4'b0000; // (3, 2) = 0
            6'b100111: o_data = 4'b0110; // (3, 3) = 6
            6'b101000: o_data = 4'b1100; // (4, 2) = 12
            6'b101001: o_data = 4'b1010; // (4, 3) = 10
            6'b101010: o_data = 4'b1011; // (5, 2) = 11
            6'b101011: o_data = 4'b0001; // (5, 3) = 1
            6'b101100: o_data = 4'b0111; // (6, 2) = 7
            6'b101101: o_data = 4'b1101; // (6, 3) = 13
            6'b101110: o_data = 4'b1101; // (7, 2) = 13
            6'b101111: o_data = 4'b1000; // (7, 3) = 8
            6'b110000: o_data = 4'b1111; // (8, 2) = 15
            6'b110001: o_data = 4'b1001; // (8, 3) = 9
            6'b110010: o_data = 4'b0001; // (9, 2) = 1
            6'b110011: o_data = 4'b0100; // (9, 3) = 4
            6'b110100: o_data = 4'b0011; // (10, 2) = 3
            6'b110101: o_data = 4'b0101; // (10, 3) = 5
            6'b110110: o_data = 4'b1110; // (11, 2) = 14
            6'b110111: o_data = 4'b1011; // (11, 3) = 11
            6'b111000: o_data = 4'b0101; // (12, 2) = 5
            6'b111001: o_data = 4'b1100; // (12, 3) = 12
            6'b111010: o_data = 4'b0010; // (13, 2) = 2
            6'b111011: o_data = 4'b0111; // (13, 3) = 7
            6'b111100: o_data = 4'b1000; // (14, 2) = 8
            6'b111101: o_data = 4'b0010; // (14, 3) = 2
            6'b111110: o_data = 4'b0100; // (15, 2) = 4
            6'b111111: o_data = 4'b1110; // (15, 3) = 14
        endcase
    end
endmodule
