magic
tech sky130A
magscale 1 2
timestamp 1639259635
<< obsli1 >>
rect 1104 1377 146803 147441
<< obsm1 >>
rect 106 1096 147278 147472
<< metal2 >>
rect 662 148803 718 149603
rect 1950 148803 2006 149603
rect 3238 148803 3294 149603
rect 4526 148803 4582 149603
rect 5814 148803 5870 149603
rect 7102 148803 7158 149603
rect 8390 148803 8446 149603
rect 9678 148803 9734 149603
rect 10966 148803 11022 149603
rect 12254 148803 12310 149603
rect 13542 148803 13598 149603
rect 14830 148803 14886 149603
rect 16118 148803 16174 149603
rect 17406 148803 17462 149603
rect 18694 148803 18750 149603
rect 19982 148803 20038 149603
rect 21270 148803 21326 149603
rect 22650 148803 22706 149603
rect 23938 148803 23994 149603
rect 25226 148803 25282 149603
rect 26514 148803 26570 149603
rect 27802 148803 27858 149603
rect 29090 148803 29146 149603
rect 30378 148803 30434 149603
rect 31666 148803 31722 149603
rect 32954 148803 33010 149603
rect 34242 148803 34298 149603
rect 35530 148803 35586 149603
rect 36818 148803 36874 149603
rect 38106 148803 38162 149603
rect 39394 148803 39450 149603
rect 40682 148803 40738 149603
rect 41970 148803 42026 149603
rect 43350 148803 43406 149603
rect 44638 148803 44694 149603
rect 45926 148803 45982 149603
rect 47214 148803 47270 149603
rect 48502 148803 48558 149603
rect 49790 148803 49846 149603
rect 51078 148803 51134 149603
rect 52366 148803 52422 149603
rect 53654 148803 53710 149603
rect 54942 148803 54998 149603
rect 56230 148803 56286 149603
rect 57518 148803 57574 149603
rect 58806 148803 58862 149603
rect 60094 148803 60150 149603
rect 61382 148803 61438 149603
rect 62670 148803 62726 149603
rect 64050 148803 64106 149603
rect 65338 148803 65394 149603
rect 66626 148803 66682 149603
rect 67914 148803 67970 149603
rect 69202 148803 69258 149603
rect 70490 148803 70546 149603
rect 71778 148803 71834 149603
rect 73066 148803 73122 149603
rect 74354 148803 74410 149603
rect 75642 148803 75698 149603
rect 76930 148803 76986 149603
rect 78218 148803 78274 149603
rect 79506 148803 79562 149603
rect 80794 148803 80850 149603
rect 82082 148803 82138 149603
rect 83370 148803 83426 149603
rect 84658 148803 84714 149603
rect 86038 148803 86094 149603
rect 87326 148803 87382 149603
rect 88614 148803 88670 149603
rect 89902 148803 89958 149603
rect 91190 148803 91246 149603
rect 92478 148803 92534 149603
rect 93766 148803 93822 149603
rect 95054 148803 95110 149603
rect 96342 148803 96398 149603
rect 97630 148803 97686 149603
rect 98918 148803 98974 149603
rect 100206 148803 100262 149603
rect 101494 148803 101550 149603
rect 102782 148803 102838 149603
rect 104070 148803 104126 149603
rect 105358 148803 105414 149603
rect 106738 148803 106794 149603
rect 108026 148803 108082 149603
rect 109314 148803 109370 149603
rect 110602 148803 110658 149603
rect 111890 148803 111946 149603
rect 113178 148803 113234 149603
rect 114466 148803 114522 149603
rect 115754 148803 115810 149603
rect 117042 148803 117098 149603
rect 118330 148803 118386 149603
rect 119618 148803 119674 149603
rect 120906 148803 120962 149603
rect 122194 148803 122250 149603
rect 123482 148803 123538 149603
rect 124770 148803 124826 149603
rect 126058 148803 126114 149603
rect 127438 148803 127494 149603
rect 128726 148803 128782 149603
rect 130014 148803 130070 149603
rect 131302 148803 131358 149603
rect 132590 148803 132646 149603
rect 133878 148803 133934 149603
rect 135166 148803 135222 149603
rect 136454 148803 136510 149603
rect 137742 148803 137798 149603
rect 139030 148803 139086 149603
rect 140318 148803 140374 149603
rect 141606 148803 141662 149603
rect 142894 148803 142950 149603
rect 144182 148803 144238 149603
rect 145470 148803 145526 149603
rect 146758 148803 146814 149603
rect 110 0 166 800
rect 386 0 442 800
rect 662 0 718 800
rect 938 0 994 800
rect 1306 0 1362 800
rect 1582 0 1638 800
rect 1858 0 1914 800
rect 2134 0 2190 800
rect 2502 0 2558 800
rect 2778 0 2834 800
rect 3054 0 3110 800
rect 3330 0 3386 800
rect 3698 0 3754 800
rect 3974 0 4030 800
rect 4250 0 4306 800
rect 4526 0 4582 800
rect 4894 0 4950 800
rect 5170 0 5226 800
rect 5446 0 5502 800
rect 5722 0 5778 800
rect 6090 0 6146 800
rect 6366 0 6422 800
rect 6642 0 6698 800
rect 6918 0 6974 800
rect 7286 0 7342 800
rect 7562 0 7618 800
rect 7838 0 7894 800
rect 8114 0 8170 800
rect 8482 0 8538 800
rect 8758 0 8814 800
rect 9034 0 9090 800
rect 9310 0 9366 800
rect 9678 0 9734 800
rect 9954 0 10010 800
rect 10230 0 10286 800
rect 10506 0 10562 800
rect 10874 0 10930 800
rect 11150 0 11206 800
rect 11426 0 11482 800
rect 11702 0 11758 800
rect 12070 0 12126 800
rect 12346 0 12402 800
rect 12622 0 12678 800
rect 12898 0 12954 800
rect 13266 0 13322 800
rect 13542 0 13598 800
rect 13818 0 13874 800
rect 14094 0 14150 800
rect 14462 0 14518 800
rect 14738 0 14794 800
rect 15014 0 15070 800
rect 15290 0 15346 800
rect 15658 0 15714 800
rect 15934 0 15990 800
rect 16210 0 16266 800
rect 16486 0 16542 800
rect 16854 0 16910 800
rect 17130 0 17186 800
rect 17406 0 17462 800
rect 17682 0 17738 800
rect 18050 0 18106 800
rect 18326 0 18382 800
rect 18602 0 18658 800
rect 18878 0 18934 800
rect 19246 0 19302 800
rect 19522 0 19578 800
rect 19798 0 19854 800
rect 20074 0 20130 800
rect 20442 0 20498 800
rect 20718 0 20774 800
rect 20994 0 21050 800
rect 21270 0 21326 800
rect 21638 0 21694 800
rect 21914 0 21970 800
rect 22190 0 22246 800
rect 22466 0 22522 800
rect 22834 0 22890 800
rect 23110 0 23166 800
rect 23386 0 23442 800
rect 23662 0 23718 800
rect 24030 0 24086 800
rect 24306 0 24362 800
rect 24582 0 24638 800
rect 24858 0 24914 800
rect 25226 0 25282 800
rect 25502 0 25558 800
rect 25778 0 25834 800
rect 26054 0 26110 800
rect 26422 0 26478 800
rect 26698 0 26754 800
rect 26974 0 27030 800
rect 27250 0 27306 800
rect 27618 0 27674 800
rect 27894 0 27950 800
rect 28170 0 28226 800
rect 28446 0 28502 800
rect 28814 0 28870 800
rect 29090 0 29146 800
rect 29366 0 29422 800
rect 29642 0 29698 800
rect 30010 0 30066 800
rect 30286 0 30342 800
rect 30562 0 30618 800
rect 30838 0 30894 800
rect 31206 0 31262 800
rect 31482 0 31538 800
rect 31758 0 31814 800
rect 32034 0 32090 800
rect 32402 0 32458 800
rect 32678 0 32734 800
rect 32954 0 33010 800
rect 33230 0 33286 800
rect 33598 0 33654 800
rect 33874 0 33930 800
rect 34150 0 34206 800
rect 34426 0 34482 800
rect 34794 0 34850 800
rect 35070 0 35126 800
rect 35346 0 35402 800
rect 35622 0 35678 800
rect 35990 0 36046 800
rect 36266 0 36322 800
rect 36542 0 36598 800
rect 36818 0 36874 800
rect 37186 0 37242 800
rect 37462 0 37518 800
rect 37738 0 37794 800
rect 38014 0 38070 800
rect 38382 0 38438 800
rect 38658 0 38714 800
rect 38934 0 38990 800
rect 39210 0 39266 800
rect 39578 0 39634 800
rect 39854 0 39910 800
rect 40130 0 40186 800
rect 40406 0 40462 800
rect 40774 0 40830 800
rect 41050 0 41106 800
rect 41326 0 41382 800
rect 41602 0 41658 800
rect 41970 0 42026 800
rect 42246 0 42302 800
rect 42522 0 42578 800
rect 42798 0 42854 800
rect 43166 0 43222 800
rect 43442 0 43498 800
rect 43718 0 43774 800
rect 43994 0 44050 800
rect 44362 0 44418 800
rect 44638 0 44694 800
rect 44914 0 44970 800
rect 45190 0 45246 800
rect 45558 0 45614 800
rect 45834 0 45890 800
rect 46110 0 46166 800
rect 46386 0 46442 800
rect 46754 0 46810 800
rect 47030 0 47086 800
rect 47306 0 47362 800
rect 47582 0 47638 800
rect 47950 0 48006 800
rect 48226 0 48282 800
rect 48502 0 48558 800
rect 48778 0 48834 800
rect 49146 0 49202 800
rect 49422 0 49478 800
rect 49698 0 49754 800
rect 50066 0 50122 800
rect 50342 0 50398 800
rect 50618 0 50674 800
rect 50894 0 50950 800
rect 51262 0 51318 800
rect 51538 0 51594 800
rect 51814 0 51870 800
rect 52090 0 52146 800
rect 52458 0 52514 800
rect 52734 0 52790 800
rect 53010 0 53066 800
rect 53286 0 53342 800
rect 53654 0 53710 800
rect 53930 0 53986 800
rect 54206 0 54262 800
rect 54482 0 54538 800
rect 54850 0 54906 800
rect 55126 0 55182 800
rect 55402 0 55458 800
rect 55678 0 55734 800
rect 56046 0 56102 800
rect 56322 0 56378 800
rect 56598 0 56654 800
rect 56874 0 56930 800
rect 57242 0 57298 800
rect 57518 0 57574 800
rect 57794 0 57850 800
rect 58070 0 58126 800
rect 58438 0 58494 800
rect 58714 0 58770 800
rect 58990 0 59046 800
rect 59266 0 59322 800
rect 59634 0 59690 800
rect 59910 0 59966 800
rect 60186 0 60242 800
rect 60462 0 60518 800
rect 60830 0 60886 800
rect 61106 0 61162 800
rect 61382 0 61438 800
rect 61658 0 61714 800
rect 62026 0 62082 800
rect 62302 0 62358 800
rect 62578 0 62634 800
rect 62854 0 62910 800
rect 63222 0 63278 800
rect 63498 0 63554 800
rect 63774 0 63830 800
rect 64050 0 64106 800
rect 64418 0 64474 800
rect 64694 0 64750 800
rect 64970 0 65026 800
rect 65246 0 65302 800
rect 65614 0 65670 800
rect 65890 0 65946 800
rect 66166 0 66222 800
rect 66442 0 66498 800
rect 66810 0 66866 800
rect 67086 0 67142 800
rect 67362 0 67418 800
rect 67638 0 67694 800
rect 68006 0 68062 800
rect 68282 0 68338 800
rect 68558 0 68614 800
rect 68834 0 68890 800
rect 69202 0 69258 800
rect 69478 0 69534 800
rect 69754 0 69810 800
rect 70030 0 70086 800
rect 70398 0 70454 800
rect 70674 0 70730 800
rect 70950 0 71006 800
rect 71226 0 71282 800
rect 71594 0 71650 800
rect 71870 0 71926 800
rect 72146 0 72202 800
rect 72422 0 72478 800
rect 72790 0 72846 800
rect 73066 0 73122 800
rect 73342 0 73398 800
rect 73618 0 73674 800
rect 73986 0 74042 800
rect 74262 0 74318 800
rect 74538 0 74594 800
rect 74814 0 74870 800
rect 75182 0 75238 800
rect 75458 0 75514 800
rect 75734 0 75790 800
rect 76010 0 76066 800
rect 76378 0 76434 800
rect 76654 0 76710 800
rect 76930 0 76986 800
rect 77206 0 77262 800
rect 77574 0 77630 800
rect 77850 0 77906 800
rect 78126 0 78182 800
rect 78402 0 78458 800
rect 78770 0 78826 800
rect 79046 0 79102 800
rect 79322 0 79378 800
rect 79598 0 79654 800
rect 79966 0 80022 800
rect 80242 0 80298 800
rect 80518 0 80574 800
rect 80794 0 80850 800
rect 81162 0 81218 800
rect 81438 0 81494 800
rect 81714 0 81770 800
rect 81990 0 82046 800
rect 82358 0 82414 800
rect 82634 0 82690 800
rect 82910 0 82966 800
rect 83186 0 83242 800
rect 83554 0 83610 800
rect 83830 0 83886 800
rect 84106 0 84162 800
rect 84382 0 84438 800
rect 84750 0 84806 800
rect 85026 0 85082 800
rect 85302 0 85358 800
rect 85578 0 85634 800
rect 85946 0 86002 800
rect 86222 0 86278 800
rect 86498 0 86554 800
rect 86774 0 86830 800
rect 87142 0 87198 800
rect 87418 0 87474 800
rect 87694 0 87750 800
rect 87970 0 88026 800
rect 88338 0 88394 800
rect 88614 0 88670 800
rect 88890 0 88946 800
rect 89166 0 89222 800
rect 89534 0 89590 800
rect 89810 0 89866 800
rect 90086 0 90142 800
rect 90362 0 90418 800
rect 90730 0 90786 800
rect 91006 0 91062 800
rect 91282 0 91338 800
rect 91558 0 91614 800
rect 91926 0 91982 800
rect 92202 0 92258 800
rect 92478 0 92534 800
rect 92754 0 92810 800
rect 93122 0 93178 800
rect 93398 0 93454 800
rect 93674 0 93730 800
rect 93950 0 94006 800
rect 94318 0 94374 800
rect 94594 0 94650 800
rect 94870 0 94926 800
rect 95146 0 95202 800
rect 95514 0 95570 800
rect 95790 0 95846 800
rect 96066 0 96122 800
rect 96342 0 96398 800
rect 96710 0 96766 800
rect 96986 0 97042 800
rect 97262 0 97318 800
rect 97538 0 97594 800
rect 97906 0 97962 800
rect 98182 0 98238 800
rect 98458 0 98514 800
rect 98826 0 98882 800
rect 99102 0 99158 800
rect 99378 0 99434 800
rect 99654 0 99710 800
rect 100022 0 100078 800
rect 100298 0 100354 800
rect 100574 0 100630 800
rect 100850 0 100906 800
rect 101218 0 101274 800
rect 101494 0 101550 800
rect 101770 0 101826 800
rect 102046 0 102102 800
rect 102414 0 102470 800
rect 102690 0 102746 800
rect 102966 0 103022 800
rect 103242 0 103298 800
rect 103610 0 103666 800
rect 103886 0 103942 800
rect 104162 0 104218 800
rect 104438 0 104494 800
rect 104806 0 104862 800
rect 105082 0 105138 800
rect 105358 0 105414 800
rect 105634 0 105690 800
rect 106002 0 106058 800
rect 106278 0 106334 800
rect 106554 0 106610 800
rect 106830 0 106886 800
rect 107198 0 107254 800
rect 107474 0 107530 800
rect 107750 0 107806 800
rect 108026 0 108082 800
rect 108394 0 108450 800
rect 108670 0 108726 800
rect 108946 0 109002 800
rect 109222 0 109278 800
rect 109590 0 109646 800
rect 109866 0 109922 800
rect 110142 0 110198 800
rect 110418 0 110474 800
rect 110786 0 110842 800
rect 111062 0 111118 800
rect 111338 0 111394 800
rect 111614 0 111670 800
rect 111982 0 112038 800
rect 112258 0 112314 800
rect 112534 0 112590 800
rect 112810 0 112866 800
rect 113178 0 113234 800
rect 113454 0 113510 800
rect 113730 0 113786 800
rect 114006 0 114062 800
rect 114374 0 114430 800
rect 114650 0 114706 800
rect 114926 0 114982 800
rect 115202 0 115258 800
rect 115570 0 115626 800
rect 115846 0 115902 800
rect 116122 0 116178 800
rect 116398 0 116454 800
rect 116766 0 116822 800
rect 117042 0 117098 800
rect 117318 0 117374 800
rect 117594 0 117650 800
rect 117962 0 118018 800
rect 118238 0 118294 800
rect 118514 0 118570 800
rect 118790 0 118846 800
rect 119158 0 119214 800
rect 119434 0 119490 800
rect 119710 0 119766 800
rect 119986 0 120042 800
rect 120354 0 120410 800
rect 120630 0 120686 800
rect 120906 0 120962 800
rect 121182 0 121238 800
rect 121550 0 121606 800
rect 121826 0 121882 800
rect 122102 0 122158 800
rect 122378 0 122434 800
rect 122746 0 122802 800
rect 123022 0 123078 800
rect 123298 0 123354 800
rect 123574 0 123630 800
rect 123942 0 123998 800
rect 124218 0 124274 800
rect 124494 0 124550 800
rect 124770 0 124826 800
rect 125138 0 125194 800
rect 125414 0 125470 800
rect 125690 0 125746 800
rect 125966 0 126022 800
rect 126334 0 126390 800
rect 126610 0 126666 800
rect 126886 0 126942 800
rect 127162 0 127218 800
rect 127530 0 127586 800
rect 127806 0 127862 800
rect 128082 0 128138 800
rect 128358 0 128414 800
rect 128726 0 128782 800
rect 129002 0 129058 800
rect 129278 0 129334 800
rect 129554 0 129610 800
rect 129922 0 129978 800
rect 130198 0 130254 800
rect 130474 0 130530 800
rect 130750 0 130806 800
rect 131118 0 131174 800
rect 131394 0 131450 800
rect 131670 0 131726 800
rect 131946 0 132002 800
rect 132314 0 132370 800
rect 132590 0 132646 800
rect 132866 0 132922 800
rect 133142 0 133198 800
rect 133510 0 133566 800
rect 133786 0 133842 800
rect 134062 0 134118 800
rect 134338 0 134394 800
rect 134706 0 134762 800
rect 134982 0 135038 800
rect 135258 0 135314 800
rect 135534 0 135590 800
rect 135902 0 135958 800
rect 136178 0 136234 800
rect 136454 0 136510 800
rect 136730 0 136786 800
rect 137098 0 137154 800
rect 137374 0 137430 800
rect 137650 0 137706 800
rect 137926 0 137982 800
rect 138294 0 138350 800
rect 138570 0 138626 800
rect 138846 0 138902 800
rect 139122 0 139178 800
rect 139490 0 139546 800
rect 139766 0 139822 800
rect 140042 0 140098 800
rect 140318 0 140374 800
rect 140686 0 140742 800
rect 140962 0 141018 800
rect 141238 0 141294 800
rect 141514 0 141570 800
rect 141882 0 141938 800
rect 142158 0 142214 800
rect 142434 0 142490 800
rect 142710 0 142766 800
rect 143078 0 143134 800
rect 143354 0 143410 800
rect 143630 0 143686 800
rect 143906 0 143962 800
rect 144274 0 144330 800
rect 144550 0 144606 800
rect 144826 0 144882 800
rect 145102 0 145158 800
rect 145470 0 145526 800
rect 145746 0 145802 800
rect 146022 0 146078 800
rect 146298 0 146354 800
rect 146666 0 146722 800
rect 146942 0 146998 800
rect 147218 0 147274 800
<< obsm2 >>
rect 112 148747 606 148866
rect 774 148747 1894 148866
rect 2062 148747 3182 148866
rect 3350 148747 4470 148866
rect 4638 148747 5758 148866
rect 5926 148747 7046 148866
rect 7214 148747 8334 148866
rect 8502 148747 9622 148866
rect 9790 148747 10910 148866
rect 11078 148747 12198 148866
rect 12366 148747 13486 148866
rect 13654 148747 14774 148866
rect 14942 148747 16062 148866
rect 16230 148747 17350 148866
rect 17518 148747 18638 148866
rect 18806 148747 19926 148866
rect 20094 148747 21214 148866
rect 21382 148747 22594 148866
rect 22762 148747 23882 148866
rect 24050 148747 25170 148866
rect 25338 148747 26458 148866
rect 26626 148747 27746 148866
rect 27914 148747 29034 148866
rect 29202 148747 30322 148866
rect 30490 148747 31610 148866
rect 31778 148747 32898 148866
rect 33066 148747 34186 148866
rect 34354 148747 35474 148866
rect 35642 148747 36762 148866
rect 36930 148747 38050 148866
rect 38218 148747 39338 148866
rect 39506 148747 40626 148866
rect 40794 148747 41914 148866
rect 42082 148747 43294 148866
rect 43462 148747 44582 148866
rect 44750 148747 45870 148866
rect 46038 148747 47158 148866
rect 47326 148747 48446 148866
rect 48614 148747 49734 148866
rect 49902 148747 51022 148866
rect 51190 148747 52310 148866
rect 52478 148747 53598 148866
rect 53766 148747 54886 148866
rect 55054 148747 56174 148866
rect 56342 148747 57462 148866
rect 57630 148747 58750 148866
rect 58918 148747 60038 148866
rect 60206 148747 61326 148866
rect 61494 148747 62614 148866
rect 62782 148747 63994 148866
rect 64162 148747 65282 148866
rect 65450 148747 66570 148866
rect 66738 148747 67858 148866
rect 68026 148747 69146 148866
rect 69314 148747 70434 148866
rect 70602 148747 71722 148866
rect 71890 148747 73010 148866
rect 73178 148747 74298 148866
rect 74466 148747 75586 148866
rect 75754 148747 76874 148866
rect 77042 148747 78162 148866
rect 78330 148747 79450 148866
rect 79618 148747 80738 148866
rect 80906 148747 82026 148866
rect 82194 148747 83314 148866
rect 83482 148747 84602 148866
rect 84770 148747 85982 148866
rect 86150 148747 87270 148866
rect 87438 148747 88558 148866
rect 88726 148747 89846 148866
rect 90014 148747 91134 148866
rect 91302 148747 92422 148866
rect 92590 148747 93710 148866
rect 93878 148747 94998 148866
rect 95166 148747 96286 148866
rect 96454 148747 97574 148866
rect 97742 148747 98862 148866
rect 99030 148747 100150 148866
rect 100318 148747 101438 148866
rect 101606 148747 102726 148866
rect 102894 148747 104014 148866
rect 104182 148747 105302 148866
rect 105470 148747 106682 148866
rect 106850 148747 107970 148866
rect 108138 148747 109258 148866
rect 109426 148747 110546 148866
rect 110714 148747 111834 148866
rect 112002 148747 113122 148866
rect 113290 148747 114410 148866
rect 114578 148747 115698 148866
rect 115866 148747 116986 148866
rect 117154 148747 118274 148866
rect 118442 148747 119562 148866
rect 119730 148747 120850 148866
rect 121018 148747 122138 148866
rect 122306 148747 123426 148866
rect 123594 148747 124714 148866
rect 124882 148747 126002 148866
rect 126170 148747 127382 148866
rect 127550 148747 128670 148866
rect 128838 148747 129958 148866
rect 130126 148747 131246 148866
rect 131414 148747 132534 148866
rect 132702 148747 133822 148866
rect 133990 148747 135110 148866
rect 135278 148747 136398 148866
rect 136566 148747 137686 148866
rect 137854 148747 138974 148866
rect 139142 148747 140262 148866
rect 140430 148747 141550 148866
rect 141718 148747 142838 148866
rect 143006 148747 144126 148866
rect 144294 148747 145414 148866
rect 145582 148747 146702 148866
rect 146870 148747 147272 148866
rect 112 856 147272 148747
rect 222 734 330 856
rect 498 734 606 856
rect 774 734 882 856
rect 1050 734 1250 856
rect 1418 734 1526 856
rect 1694 734 1802 856
rect 1970 734 2078 856
rect 2246 734 2446 856
rect 2614 734 2722 856
rect 2890 734 2998 856
rect 3166 734 3274 856
rect 3442 734 3642 856
rect 3810 734 3918 856
rect 4086 734 4194 856
rect 4362 734 4470 856
rect 4638 734 4838 856
rect 5006 734 5114 856
rect 5282 734 5390 856
rect 5558 734 5666 856
rect 5834 734 6034 856
rect 6202 734 6310 856
rect 6478 734 6586 856
rect 6754 734 6862 856
rect 7030 734 7230 856
rect 7398 734 7506 856
rect 7674 734 7782 856
rect 7950 734 8058 856
rect 8226 734 8426 856
rect 8594 734 8702 856
rect 8870 734 8978 856
rect 9146 734 9254 856
rect 9422 734 9622 856
rect 9790 734 9898 856
rect 10066 734 10174 856
rect 10342 734 10450 856
rect 10618 734 10818 856
rect 10986 734 11094 856
rect 11262 734 11370 856
rect 11538 734 11646 856
rect 11814 734 12014 856
rect 12182 734 12290 856
rect 12458 734 12566 856
rect 12734 734 12842 856
rect 13010 734 13210 856
rect 13378 734 13486 856
rect 13654 734 13762 856
rect 13930 734 14038 856
rect 14206 734 14406 856
rect 14574 734 14682 856
rect 14850 734 14958 856
rect 15126 734 15234 856
rect 15402 734 15602 856
rect 15770 734 15878 856
rect 16046 734 16154 856
rect 16322 734 16430 856
rect 16598 734 16798 856
rect 16966 734 17074 856
rect 17242 734 17350 856
rect 17518 734 17626 856
rect 17794 734 17994 856
rect 18162 734 18270 856
rect 18438 734 18546 856
rect 18714 734 18822 856
rect 18990 734 19190 856
rect 19358 734 19466 856
rect 19634 734 19742 856
rect 19910 734 20018 856
rect 20186 734 20386 856
rect 20554 734 20662 856
rect 20830 734 20938 856
rect 21106 734 21214 856
rect 21382 734 21582 856
rect 21750 734 21858 856
rect 22026 734 22134 856
rect 22302 734 22410 856
rect 22578 734 22778 856
rect 22946 734 23054 856
rect 23222 734 23330 856
rect 23498 734 23606 856
rect 23774 734 23974 856
rect 24142 734 24250 856
rect 24418 734 24526 856
rect 24694 734 24802 856
rect 24970 734 25170 856
rect 25338 734 25446 856
rect 25614 734 25722 856
rect 25890 734 25998 856
rect 26166 734 26366 856
rect 26534 734 26642 856
rect 26810 734 26918 856
rect 27086 734 27194 856
rect 27362 734 27562 856
rect 27730 734 27838 856
rect 28006 734 28114 856
rect 28282 734 28390 856
rect 28558 734 28758 856
rect 28926 734 29034 856
rect 29202 734 29310 856
rect 29478 734 29586 856
rect 29754 734 29954 856
rect 30122 734 30230 856
rect 30398 734 30506 856
rect 30674 734 30782 856
rect 30950 734 31150 856
rect 31318 734 31426 856
rect 31594 734 31702 856
rect 31870 734 31978 856
rect 32146 734 32346 856
rect 32514 734 32622 856
rect 32790 734 32898 856
rect 33066 734 33174 856
rect 33342 734 33542 856
rect 33710 734 33818 856
rect 33986 734 34094 856
rect 34262 734 34370 856
rect 34538 734 34738 856
rect 34906 734 35014 856
rect 35182 734 35290 856
rect 35458 734 35566 856
rect 35734 734 35934 856
rect 36102 734 36210 856
rect 36378 734 36486 856
rect 36654 734 36762 856
rect 36930 734 37130 856
rect 37298 734 37406 856
rect 37574 734 37682 856
rect 37850 734 37958 856
rect 38126 734 38326 856
rect 38494 734 38602 856
rect 38770 734 38878 856
rect 39046 734 39154 856
rect 39322 734 39522 856
rect 39690 734 39798 856
rect 39966 734 40074 856
rect 40242 734 40350 856
rect 40518 734 40718 856
rect 40886 734 40994 856
rect 41162 734 41270 856
rect 41438 734 41546 856
rect 41714 734 41914 856
rect 42082 734 42190 856
rect 42358 734 42466 856
rect 42634 734 42742 856
rect 42910 734 43110 856
rect 43278 734 43386 856
rect 43554 734 43662 856
rect 43830 734 43938 856
rect 44106 734 44306 856
rect 44474 734 44582 856
rect 44750 734 44858 856
rect 45026 734 45134 856
rect 45302 734 45502 856
rect 45670 734 45778 856
rect 45946 734 46054 856
rect 46222 734 46330 856
rect 46498 734 46698 856
rect 46866 734 46974 856
rect 47142 734 47250 856
rect 47418 734 47526 856
rect 47694 734 47894 856
rect 48062 734 48170 856
rect 48338 734 48446 856
rect 48614 734 48722 856
rect 48890 734 49090 856
rect 49258 734 49366 856
rect 49534 734 49642 856
rect 49810 734 50010 856
rect 50178 734 50286 856
rect 50454 734 50562 856
rect 50730 734 50838 856
rect 51006 734 51206 856
rect 51374 734 51482 856
rect 51650 734 51758 856
rect 51926 734 52034 856
rect 52202 734 52402 856
rect 52570 734 52678 856
rect 52846 734 52954 856
rect 53122 734 53230 856
rect 53398 734 53598 856
rect 53766 734 53874 856
rect 54042 734 54150 856
rect 54318 734 54426 856
rect 54594 734 54794 856
rect 54962 734 55070 856
rect 55238 734 55346 856
rect 55514 734 55622 856
rect 55790 734 55990 856
rect 56158 734 56266 856
rect 56434 734 56542 856
rect 56710 734 56818 856
rect 56986 734 57186 856
rect 57354 734 57462 856
rect 57630 734 57738 856
rect 57906 734 58014 856
rect 58182 734 58382 856
rect 58550 734 58658 856
rect 58826 734 58934 856
rect 59102 734 59210 856
rect 59378 734 59578 856
rect 59746 734 59854 856
rect 60022 734 60130 856
rect 60298 734 60406 856
rect 60574 734 60774 856
rect 60942 734 61050 856
rect 61218 734 61326 856
rect 61494 734 61602 856
rect 61770 734 61970 856
rect 62138 734 62246 856
rect 62414 734 62522 856
rect 62690 734 62798 856
rect 62966 734 63166 856
rect 63334 734 63442 856
rect 63610 734 63718 856
rect 63886 734 63994 856
rect 64162 734 64362 856
rect 64530 734 64638 856
rect 64806 734 64914 856
rect 65082 734 65190 856
rect 65358 734 65558 856
rect 65726 734 65834 856
rect 66002 734 66110 856
rect 66278 734 66386 856
rect 66554 734 66754 856
rect 66922 734 67030 856
rect 67198 734 67306 856
rect 67474 734 67582 856
rect 67750 734 67950 856
rect 68118 734 68226 856
rect 68394 734 68502 856
rect 68670 734 68778 856
rect 68946 734 69146 856
rect 69314 734 69422 856
rect 69590 734 69698 856
rect 69866 734 69974 856
rect 70142 734 70342 856
rect 70510 734 70618 856
rect 70786 734 70894 856
rect 71062 734 71170 856
rect 71338 734 71538 856
rect 71706 734 71814 856
rect 71982 734 72090 856
rect 72258 734 72366 856
rect 72534 734 72734 856
rect 72902 734 73010 856
rect 73178 734 73286 856
rect 73454 734 73562 856
rect 73730 734 73930 856
rect 74098 734 74206 856
rect 74374 734 74482 856
rect 74650 734 74758 856
rect 74926 734 75126 856
rect 75294 734 75402 856
rect 75570 734 75678 856
rect 75846 734 75954 856
rect 76122 734 76322 856
rect 76490 734 76598 856
rect 76766 734 76874 856
rect 77042 734 77150 856
rect 77318 734 77518 856
rect 77686 734 77794 856
rect 77962 734 78070 856
rect 78238 734 78346 856
rect 78514 734 78714 856
rect 78882 734 78990 856
rect 79158 734 79266 856
rect 79434 734 79542 856
rect 79710 734 79910 856
rect 80078 734 80186 856
rect 80354 734 80462 856
rect 80630 734 80738 856
rect 80906 734 81106 856
rect 81274 734 81382 856
rect 81550 734 81658 856
rect 81826 734 81934 856
rect 82102 734 82302 856
rect 82470 734 82578 856
rect 82746 734 82854 856
rect 83022 734 83130 856
rect 83298 734 83498 856
rect 83666 734 83774 856
rect 83942 734 84050 856
rect 84218 734 84326 856
rect 84494 734 84694 856
rect 84862 734 84970 856
rect 85138 734 85246 856
rect 85414 734 85522 856
rect 85690 734 85890 856
rect 86058 734 86166 856
rect 86334 734 86442 856
rect 86610 734 86718 856
rect 86886 734 87086 856
rect 87254 734 87362 856
rect 87530 734 87638 856
rect 87806 734 87914 856
rect 88082 734 88282 856
rect 88450 734 88558 856
rect 88726 734 88834 856
rect 89002 734 89110 856
rect 89278 734 89478 856
rect 89646 734 89754 856
rect 89922 734 90030 856
rect 90198 734 90306 856
rect 90474 734 90674 856
rect 90842 734 90950 856
rect 91118 734 91226 856
rect 91394 734 91502 856
rect 91670 734 91870 856
rect 92038 734 92146 856
rect 92314 734 92422 856
rect 92590 734 92698 856
rect 92866 734 93066 856
rect 93234 734 93342 856
rect 93510 734 93618 856
rect 93786 734 93894 856
rect 94062 734 94262 856
rect 94430 734 94538 856
rect 94706 734 94814 856
rect 94982 734 95090 856
rect 95258 734 95458 856
rect 95626 734 95734 856
rect 95902 734 96010 856
rect 96178 734 96286 856
rect 96454 734 96654 856
rect 96822 734 96930 856
rect 97098 734 97206 856
rect 97374 734 97482 856
rect 97650 734 97850 856
rect 98018 734 98126 856
rect 98294 734 98402 856
rect 98570 734 98770 856
rect 98938 734 99046 856
rect 99214 734 99322 856
rect 99490 734 99598 856
rect 99766 734 99966 856
rect 100134 734 100242 856
rect 100410 734 100518 856
rect 100686 734 100794 856
rect 100962 734 101162 856
rect 101330 734 101438 856
rect 101606 734 101714 856
rect 101882 734 101990 856
rect 102158 734 102358 856
rect 102526 734 102634 856
rect 102802 734 102910 856
rect 103078 734 103186 856
rect 103354 734 103554 856
rect 103722 734 103830 856
rect 103998 734 104106 856
rect 104274 734 104382 856
rect 104550 734 104750 856
rect 104918 734 105026 856
rect 105194 734 105302 856
rect 105470 734 105578 856
rect 105746 734 105946 856
rect 106114 734 106222 856
rect 106390 734 106498 856
rect 106666 734 106774 856
rect 106942 734 107142 856
rect 107310 734 107418 856
rect 107586 734 107694 856
rect 107862 734 107970 856
rect 108138 734 108338 856
rect 108506 734 108614 856
rect 108782 734 108890 856
rect 109058 734 109166 856
rect 109334 734 109534 856
rect 109702 734 109810 856
rect 109978 734 110086 856
rect 110254 734 110362 856
rect 110530 734 110730 856
rect 110898 734 111006 856
rect 111174 734 111282 856
rect 111450 734 111558 856
rect 111726 734 111926 856
rect 112094 734 112202 856
rect 112370 734 112478 856
rect 112646 734 112754 856
rect 112922 734 113122 856
rect 113290 734 113398 856
rect 113566 734 113674 856
rect 113842 734 113950 856
rect 114118 734 114318 856
rect 114486 734 114594 856
rect 114762 734 114870 856
rect 115038 734 115146 856
rect 115314 734 115514 856
rect 115682 734 115790 856
rect 115958 734 116066 856
rect 116234 734 116342 856
rect 116510 734 116710 856
rect 116878 734 116986 856
rect 117154 734 117262 856
rect 117430 734 117538 856
rect 117706 734 117906 856
rect 118074 734 118182 856
rect 118350 734 118458 856
rect 118626 734 118734 856
rect 118902 734 119102 856
rect 119270 734 119378 856
rect 119546 734 119654 856
rect 119822 734 119930 856
rect 120098 734 120298 856
rect 120466 734 120574 856
rect 120742 734 120850 856
rect 121018 734 121126 856
rect 121294 734 121494 856
rect 121662 734 121770 856
rect 121938 734 122046 856
rect 122214 734 122322 856
rect 122490 734 122690 856
rect 122858 734 122966 856
rect 123134 734 123242 856
rect 123410 734 123518 856
rect 123686 734 123886 856
rect 124054 734 124162 856
rect 124330 734 124438 856
rect 124606 734 124714 856
rect 124882 734 125082 856
rect 125250 734 125358 856
rect 125526 734 125634 856
rect 125802 734 125910 856
rect 126078 734 126278 856
rect 126446 734 126554 856
rect 126722 734 126830 856
rect 126998 734 127106 856
rect 127274 734 127474 856
rect 127642 734 127750 856
rect 127918 734 128026 856
rect 128194 734 128302 856
rect 128470 734 128670 856
rect 128838 734 128946 856
rect 129114 734 129222 856
rect 129390 734 129498 856
rect 129666 734 129866 856
rect 130034 734 130142 856
rect 130310 734 130418 856
rect 130586 734 130694 856
rect 130862 734 131062 856
rect 131230 734 131338 856
rect 131506 734 131614 856
rect 131782 734 131890 856
rect 132058 734 132258 856
rect 132426 734 132534 856
rect 132702 734 132810 856
rect 132978 734 133086 856
rect 133254 734 133454 856
rect 133622 734 133730 856
rect 133898 734 134006 856
rect 134174 734 134282 856
rect 134450 734 134650 856
rect 134818 734 134926 856
rect 135094 734 135202 856
rect 135370 734 135478 856
rect 135646 734 135846 856
rect 136014 734 136122 856
rect 136290 734 136398 856
rect 136566 734 136674 856
rect 136842 734 137042 856
rect 137210 734 137318 856
rect 137486 734 137594 856
rect 137762 734 137870 856
rect 138038 734 138238 856
rect 138406 734 138514 856
rect 138682 734 138790 856
rect 138958 734 139066 856
rect 139234 734 139434 856
rect 139602 734 139710 856
rect 139878 734 139986 856
rect 140154 734 140262 856
rect 140430 734 140630 856
rect 140798 734 140906 856
rect 141074 734 141182 856
rect 141350 734 141458 856
rect 141626 734 141826 856
rect 141994 734 142102 856
rect 142270 734 142378 856
rect 142546 734 142654 856
rect 142822 734 143022 856
rect 143190 734 143298 856
rect 143466 734 143574 856
rect 143742 734 143850 856
rect 144018 734 144218 856
rect 144386 734 144494 856
rect 144662 734 144770 856
rect 144938 734 145046 856
rect 145214 734 145414 856
rect 145582 734 145690 856
rect 145858 734 145966 856
rect 146134 734 146242 856
rect 146410 734 146610 856
rect 146778 734 146886 856
rect 147054 734 147162 856
<< obsm3 >>
rect 841 1803 144703 147457
<< metal4 >>
rect 4208 2128 4528 147472
rect 19568 2128 19888 147472
rect 34928 2128 35248 147472
rect 50288 2128 50608 147472
rect 65648 2128 65968 147472
rect 81008 2128 81328 147472
rect 96368 2128 96688 147472
rect 111728 2128 112048 147472
rect 127088 2128 127408 147472
rect 142448 2128 142768 147472
<< obsm4 >>
rect 4659 3571 19488 104141
rect 19968 3571 34848 104141
rect 35328 3571 50208 104141
rect 50688 3571 65568 104141
rect 66048 3571 80928 104141
rect 81408 3571 96288 104141
rect 96768 3571 111648 104141
rect 112128 3571 127008 104141
rect 127488 3571 135549 104141
<< labels >>
rlabel metal2 s 662 148803 718 149603 6 io_in[0]
port 1 nsew signal input
rlabel metal2 s 39394 148803 39450 149603 6 io_in[10]
port 2 nsew signal input
rlabel metal2 s 43350 148803 43406 149603 6 io_in[11]
port 3 nsew signal input
rlabel metal2 s 47214 148803 47270 149603 6 io_in[12]
port 4 nsew signal input
rlabel metal2 s 51078 148803 51134 149603 6 io_in[13]
port 5 nsew signal input
rlabel metal2 s 54942 148803 54998 149603 6 io_in[14]
port 6 nsew signal input
rlabel metal2 s 58806 148803 58862 149603 6 io_in[15]
port 7 nsew signal input
rlabel metal2 s 62670 148803 62726 149603 6 io_in[16]
port 8 nsew signal input
rlabel metal2 s 66626 148803 66682 149603 6 io_in[17]
port 9 nsew signal input
rlabel metal2 s 70490 148803 70546 149603 6 io_in[18]
port 10 nsew signal input
rlabel metal2 s 74354 148803 74410 149603 6 io_in[19]
port 11 nsew signal input
rlabel metal2 s 4526 148803 4582 149603 6 io_in[1]
port 12 nsew signal input
rlabel metal2 s 78218 148803 78274 149603 6 io_in[20]
port 13 nsew signal input
rlabel metal2 s 82082 148803 82138 149603 6 io_in[21]
port 14 nsew signal input
rlabel metal2 s 86038 148803 86094 149603 6 io_in[22]
port 15 nsew signal input
rlabel metal2 s 89902 148803 89958 149603 6 io_in[23]
port 16 nsew signal input
rlabel metal2 s 93766 148803 93822 149603 6 io_in[24]
port 17 nsew signal input
rlabel metal2 s 97630 148803 97686 149603 6 io_in[25]
port 18 nsew signal input
rlabel metal2 s 101494 148803 101550 149603 6 io_in[26]
port 19 nsew signal input
rlabel metal2 s 105358 148803 105414 149603 6 io_in[27]
port 20 nsew signal input
rlabel metal2 s 109314 148803 109370 149603 6 io_in[28]
port 21 nsew signal input
rlabel metal2 s 113178 148803 113234 149603 6 io_in[29]
port 22 nsew signal input
rlabel metal2 s 8390 148803 8446 149603 6 io_in[2]
port 23 nsew signal input
rlabel metal2 s 117042 148803 117098 149603 6 io_in[30]
port 24 nsew signal input
rlabel metal2 s 120906 148803 120962 149603 6 io_in[31]
port 25 nsew signal input
rlabel metal2 s 124770 148803 124826 149603 6 io_in[32]
port 26 nsew signal input
rlabel metal2 s 128726 148803 128782 149603 6 io_in[33]
port 27 nsew signal input
rlabel metal2 s 132590 148803 132646 149603 6 io_in[34]
port 28 nsew signal input
rlabel metal2 s 136454 148803 136510 149603 6 io_in[35]
port 29 nsew signal input
rlabel metal2 s 140318 148803 140374 149603 6 io_in[36]
port 30 nsew signal input
rlabel metal2 s 144182 148803 144238 149603 6 io_in[37]
port 31 nsew signal input
rlabel metal2 s 12254 148803 12310 149603 6 io_in[3]
port 32 nsew signal input
rlabel metal2 s 16118 148803 16174 149603 6 io_in[4]
port 33 nsew signal input
rlabel metal2 s 19982 148803 20038 149603 6 io_in[5]
port 34 nsew signal input
rlabel metal2 s 23938 148803 23994 149603 6 io_in[6]
port 35 nsew signal input
rlabel metal2 s 27802 148803 27858 149603 6 io_in[7]
port 36 nsew signal input
rlabel metal2 s 31666 148803 31722 149603 6 io_in[8]
port 37 nsew signal input
rlabel metal2 s 35530 148803 35586 149603 6 io_in[9]
port 38 nsew signal input
rlabel metal2 s 1950 148803 2006 149603 6 io_oeb[0]
port 39 nsew signal output
rlabel metal2 s 40682 148803 40738 149603 6 io_oeb[10]
port 40 nsew signal output
rlabel metal2 s 44638 148803 44694 149603 6 io_oeb[11]
port 41 nsew signal output
rlabel metal2 s 48502 148803 48558 149603 6 io_oeb[12]
port 42 nsew signal output
rlabel metal2 s 52366 148803 52422 149603 6 io_oeb[13]
port 43 nsew signal output
rlabel metal2 s 56230 148803 56286 149603 6 io_oeb[14]
port 44 nsew signal output
rlabel metal2 s 60094 148803 60150 149603 6 io_oeb[15]
port 45 nsew signal output
rlabel metal2 s 64050 148803 64106 149603 6 io_oeb[16]
port 46 nsew signal output
rlabel metal2 s 67914 148803 67970 149603 6 io_oeb[17]
port 47 nsew signal output
rlabel metal2 s 71778 148803 71834 149603 6 io_oeb[18]
port 48 nsew signal output
rlabel metal2 s 75642 148803 75698 149603 6 io_oeb[19]
port 49 nsew signal output
rlabel metal2 s 5814 148803 5870 149603 6 io_oeb[1]
port 50 nsew signal output
rlabel metal2 s 79506 148803 79562 149603 6 io_oeb[20]
port 51 nsew signal output
rlabel metal2 s 83370 148803 83426 149603 6 io_oeb[21]
port 52 nsew signal output
rlabel metal2 s 87326 148803 87382 149603 6 io_oeb[22]
port 53 nsew signal output
rlabel metal2 s 91190 148803 91246 149603 6 io_oeb[23]
port 54 nsew signal output
rlabel metal2 s 95054 148803 95110 149603 6 io_oeb[24]
port 55 nsew signal output
rlabel metal2 s 98918 148803 98974 149603 6 io_oeb[25]
port 56 nsew signal output
rlabel metal2 s 102782 148803 102838 149603 6 io_oeb[26]
port 57 nsew signal output
rlabel metal2 s 106738 148803 106794 149603 6 io_oeb[27]
port 58 nsew signal output
rlabel metal2 s 110602 148803 110658 149603 6 io_oeb[28]
port 59 nsew signal output
rlabel metal2 s 114466 148803 114522 149603 6 io_oeb[29]
port 60 nsew signal output
rlabel metal2 s 9678 148803 9734 149603 6 io_oeb[2]
port 61 nsew signal output
rlabel metal2 s 118330 148803 118386 149603 6 io_oeb[30]
port 62 nsew signal output
rlabel metal2 s 122194 148803 122250 149603 6 io_oeb[31]
port 63 nsew signal output
rlabel metal2 s 126058 148803 126114 149603 6 io_oeb[32]
port 64 nsew signal output
rlabel metal2 s 130014 148803 130070 149603 6 io_oeb[33]
port 65 nsew signal output
rlabel metal2 s 133878 148803 133934 149603 6 io_oeb[34]
port 66 nsew signal output
rlabel metal2 s 137742 148803 137798 149603 6 io_oeb[35]
port 67 nsew signal output
rlabel metal2 s 141606 148803 141662 149603 6 io_oeb[36]
port 68 nsew signal output
rlabel metal2 s 145470 148803 145526 149603 6 io_oeb[37]
port 69 nsew signal output
rlabel metal2 s 13542 148803 13598 149603 6 io_oeb[3]
port 70 nsew signal output
rlabel metal2 s 17406 148803 17462 149603 6 io_oeb[4]
port 71 nsew signal output
rlabel metal2 s 21270 148803 21326 149603 6 io_oeb[5]
port 72 nsew signal output
rlabel metal2 s 25226 148803 25282 149603 6 io_oeb[6]
port 73 nsew signal output
rlabel metal2 s 29090 148803 29146 149603 6 io_oeb[7]
port 74 nsew signal output
rlabel metal2 s 32954 148803 33010 149603 6 io_oeb[8]
port 75 nsew signal output
rlabel metal2 s 36818 148803 36874 149603 6 io_oeb[9]
port 76 nsew signal output
rlabel metal2 s 3238 148803 3294 149603 6 io_out[0]
port 77 nsew signal output
rlabel metal2 s 41970 148803 42026 149603 6 io_out[10]
port 78 nsew signal output
rlabel metal2 s 45926 148803 45982 149603 6 io_out[11]
port 79 nsew signal output
rlabel metal2 s 49790 148803 49846 149603 6 io_out[12]
port 80 nsew signal output
rlabel metal2 s 53654 148803 53710 149603 6 io_out[13]
port 81 nsew signal output
rlabel metal2 s 57518 148803 57574 149603 6 io_out[14]
port 82 nsew signal output
rlabel metal2 s 61382 148803 61438 149603 6 io_out[15]
port 83 nsew signal output
rlabel metal2 s 65338 148803 65394 149603 6 io_out[16]
port 84 nsew signal output
rlabel metal2 s 69202 148803 69258 149603 6 io_out[17]
port 85 nsew signal output
rlabel metal2 s 73066 148803 73122 149603 6 io_out[18]
port 86 nsew signal output
rlabel metal2 s 76930 148803 76986 149603 6 io_out[19]
port 87 nsew signal output
rlabel metal2 s 7102 148803 7158 149603 6 io_out[1]
port 88 nsew signal output
rlabel metal2 s 80794 148803 80850 149603 6 io_out[20]
port 89 nsew signal output
rlabel metal2 s 84658 148803 84714 149603 6 io_out[21]
port 90 nsew signal output
rlabel metal2 s 88614 148803 88670 149603 6 io_out[22]
port 91 nsew signal output
rlabel metal2 s 92478 148803 92534 149603 6 io_out[23]
port 92 nsew signal output
rlabel metal2 s 96342 148803 96398 149603 6 io_out[24]
port 93 nsew signal output
rlabel metal2 s 100206 148803 100262 149603 6 io_out[25]
port 94 nsew signal output
rlabel metal2 s 104070 148803 104126 149603 6 io_out[26]
port 95 nsew signal output
rlabel metal2 s 108026 148803 108082 149603 6 io_out[27]
port 96 nsew signal output
rlabel metal2 s 111890 148803 111946 149603 6 io_out[28]
port 97 nsew signal output
rlabel metal2 s 115754 148803 115810 149603 6 io_out[29]
port 98 nsew signal output
rlabel metal2 s 10966 148803 11022 149603 6 io_out[2]
port 99 nsew signal output
rlabel metal2 s 119618 148803 119674 149603 6 io_out[30]
port 100 nsew signal output
rlabel metal2 s 123482 148803 123538 149603 6 io_out[31]
port 101 nsew signal output
rlabel metal2 s 127438 148803 127494 149603 6 io_out[32]
port 102 nsew signal output
rlabel metal2 s 131302 148803 131358 149603 6 io_out[33]
port 103 nsew signal output
rlabel metal2 s 135166 148803 135222 149603 6 io_out[34]
port 104 nsew signal output
rlabel metal2 s 139030 148803 139086 149603 6 io_out[35]
port 105 nsew signal output
rlabel metal2 s 142894 148803 142950 149603 6 io_out[36]
port 106 nsew signal output
rlabel metal2 s 146758 148803 146814 149603 6 io_out[37]
port 107 nsew signal output
rlabel metal2 s 14830 148803 14886 149603 6 io_out[3]
port 108 nsew signal output
rlabel metal2 s 18694 148803 18750 149603 6 io_out[4]
port 109 nsew signal output
rlabel metal2 s 22650 148803 22706 149603 6 io_out[5]
port 110 nsew signal output
rlabel metal2 s 26514 148803 26570 149603 6 io_out[6]
port 111 nsew signal output
rlabel metal2 s 30378 148803 30434 149603 6 io_out[7]
port 112 nsew signal output
rlabel metal2 s 34242 148803 34298 149603 6 io_out[8]
port 113 nsew signal output
rlabel metal2 s 38106 148803 38162 149603 6 io_out[9]
port 114 nsew signal output
rlabel metal2 s 146666 0 146722 800 6 irq[0]
port 115 nsew signal output
rlabel metal2 s 146942 0 146998 800 6 irq[1]
port 116 nsew signal output
rlabel metal2 s 147218 0 147274 800 6 irq[2]
port 117 nsew signal output
rlabel metal2 s 31758 0 31814 800 6 la_data_in[0]
port 118 nsew signal input
rlabel metal2 s 121550 0 121606 800 6 la_data_in[100]
port 119 nsew signal input
rlabel metal2 s 122378 0 122434 800 6 la_data_in[101]
port 120 nsew signal input
rlabel metal2 s 123298 0 123354 800 6 la_data_in[102]
port 121 nsew signal input
rlabel metal2 s 124218 0 124274 800 6 la_data_in[103]
port 122 nsew signal input
rlabel metal2 s 125138 0 125194 800 6 la_data_in[104]
port 123 nsew signal input
rlabel metal2 s 125966 0 126022 800 6 la_data_in[105]
port 124 nsew signal input
rlabel metal2 s 126886 0 126942 800 6 la_data_in[106]
port 125 nsew signal input
rlabel metal2 s 127806 0 127862 800 6 la_data_in[107]
port 126 nsew signal input
rlabel metal2 s 128726 0 128782 800 6 la_data_in[108]
port 127 nsew signal input
rlabel metal2 s 129554 0 129610 800 6 la_data_in[109]
port 128 nsew signal input
rlabel metal2 s 40774 0 40830 800 6 la_data_in[10]
port 129 nsew signal input
rlabel metal2 s 130474 0 130530 800 6 la_data_in[110]
port 130 nsew signal input
rlabel metal2 s 131394 0 131450 800 6 la_data_in[111]
port 131 nsew signal input
rlabel metal2 s 132314 0 132370 800 6 la_data_in[112]
port 132 nsew signal input
rlabel metal2 s 133142 0 133198 800 6 la_data_in[113]
port 133 nsew signal input
rlabel metal2 s 134062 0 134118 800 6 la_data_in[114]
port 134 nsew signal input
rlabel metal2 s 134982 0 135038 800 6 la_data_in[115]
port 135 nsew signal input
rlabel metal2 s 135902 0 135958 800 6 la_data_in[116]
port 136 nsew signal input
rlabel metal2 s 136730 0 136786 800 6 la_data_in[117]
port 137 nsew signal input
rlabel metal2 s 137650 0 137706 800 6 la_data_in[118]
port 138 nsew signal input
rlabel metal2 s 138570 0 138626 800 6 la_data_in[119]
port 139 nsew signal input
rlabel metal2 s 41602 0 41658 800 6 la_data_in[11]
port 140 nsew signal input
rlabel metal2 s 139490 0 139546 800 6 la_data_in[120]
port 141 nsew signal input
rlabel metal2 s 140318 0 140374 800 6 la_data_in[121]
port 142 nsew signal input
rlabel metal2 s 141238 0 141294 800 6 la_data_in[122]
port 143 nsew signal input
rlabel metal2 s 142158 0 142214 800 6 la_data_in[123]
port 144 nsew signal input
rlabel metal2 s 143078 0 143134 800 6 la_data_in[124]
port 145 nsew signal input
rlabel metal2 s 143906 0 143962 800 6 la_data_in[125]
port 146 nsew signal input
rlabel metal2 s 144826 0 144882 800 6 la_data_in[126]
port 147 nsew signal input
rlabel metal2 s 145746 0 145802 800 6 la_data_in[127]
port 148 nsew signal input
rlabel metal2 s 42522 0 42578 800 6 la_data_in[12]
port 149 nsew signal input
rlabel metal2 s 43442 0 43498 800 6 la_data_in[13]
port 150 nsew signal input
rlabel metal2 s 44362 0 44418 800 6 la_data_in[14]
port 151 nsew signal input
rlabel metal2 s 45190 0 45246 800 6 la_data_in[15]
port 152 nsew signal input
rlabel metal2 s 46110 0 46166 800 6 la_data_in[16]
port 153 nsew signal input
rlabel metal2 s 47030 0 47086 800 6 la_data_in[17]
port 154 nsew signal input
rlabel metal2 s 47950 0 48006 800 6 la_data_in[18]
port 155 nsew signal input
rlabel metal2 s 48778 0 48834 800 6 la_data_in[19]
port 156 nsew signal input
rlabel metal2 s 32678 0 32734 800 6 la_data_in[1]
port 157 nsew signal input
rlabel metal2 s 49698 0 49754 800 6 la_data_in[20]
port 158 nsew signal input
rlabel metal2 s 50618 0 50674 800 6 la_data_in[21]
port 159 nsew signal input
rlabel metal2 s 51538 0 51594 800 6 la_data_in[22]
port 160 nsew signal input
rlabel metal2 s 52458 0 52514 800 6 la_data_in[23]
port 161 nsew signal input
rlabel metal2 s 53286 0 53342 800 6 la_data_in[24]
port 162 nsew signal input
rlabel metal2 s 54206 0 54262 800 6 la_data_in[25]
port 163 nsew signal input
rlabel metal2 s 55126 0 55182 800 6 la_data_in[26]
port 164 nsew signal input
rlabel metal2 s 56046 0 56102 800 6 la_data_in[27]
port 165 nsew signal input
rlabel metal2 s 56874 0 56930 800 6 la_data_in[28]
port 166 nsew signal input
rlabel metal2 s 57794 0 57850 800 6 la_data_in[29]
port 167 nsew signal input
rlabel metal2 s 33598 0 33654 800 6 la_data_in[2]
port 168 nsew signal input
rlabel metal2 s 58714 0 58770 800 6 la_data_in[30]
port 169 nsew signal input
rlabel metal2 s 59634 0 59690 800 6 la_data_in[31]
port 170 nsew signal input
rlabel metal2 s 60462 0 60518 800 6 la_data_in[32]
port 171 nsew signal input
rlabel metal2 s 61382 0 61438 800 6 la_data_in[33]
port 172 nsew signal input
rlabel metal2 s 62302 0 62358 800 6 la_data_in[34]
port 173 nsew signal input
rlabel metal2 s 63222 0 63278 800 6 la_data_in[35]
port 174 nsew signal input
rlabel metal2 s 64050 0 64106 800 6 la_data_in[36]
port 175 nsew signal input
rlabel metal2 s 64970 0 65026 800 6 la_data_in[37]
port 176 nsew signal input
rlabel metal2 s 65890 0 65946 800 6 la_data_in[38]
port 177 nsew signal input
rlabel metal2 s 66810 0 66866 800 6 la_data_in[39]
port 178 nsew signal input
rlabel metal2 s 34426 0 34482 800 6 la_data_in[3]
port 179 nsew signal input
rlabel metal2 s 67638 0 67694 800 6 la_data_in[40]
port 180 nsew signal input
rlabel metal2 s 68558 0 68614 800 6 la_data_in[41]
port 181 nsew signal input
rlabel metal2 s 69478 0 69534 800 6 la_data_in[42]
port 182 nsew signal input
rlabel metal2 s 70398 0 70454 800 6 la_data_in[43]
port 183 nsew signal input
rlabel metal2 s 71226 0 71282 800 6 la_data_in[44]
port 184 nsew signal input
rlabel metal2 s 72146 0 72202 800 6 la_data_in[45]
port 185 nsew signal input
rlabel metal2 s 73066 0 73122 800 6 la_data_in[46]
port 186 nsew signal input
rlabel metal2 s 73986 0 74042 800 6 la_data_in[47]
port 187 nsew signal input
rlabel metal2 s 74814 0 74870 800 6 la_data_in[48]
port 188 nsew signal input
rlabel metal2 s 75734 0 75790 800 6 la_data_in[49]
port 189 nsew signal input
rlabel metal2 s 35346 0 35402 800 6 la_data_in[4]
port 190 nsew signal input
rlabel metal2 s 76654 0 76710 800 6 la_data_in[50]
port 191 nsew signal input
rlabel metal2 s 77574 0 77630 800 6 la_data_in[51]
port 192 nsew signal input
rlabel metal2 s 78402 0 78458 800 6 la_data_in[52]
port 193 nsew signal input
rlabel metal2 s 79322 0 79378 800 6 la_data_in[53]
port 194 nsew signal input
rlabel metal2 s 80242 0 80298 800 6 la_data_in[54]
port 195 nsew signal input
rlabel metal2 s 81162 0 81218 800 6 la_data_in[55]
port 196 nsew signal input
rlabel metal2 s 81990 0 82046 800 6 la_data_in[56]
port 197 nsew signal input
rlabel metal2 s 82910 0 82966 800 6 la_data_in[57]
port 198 nsew signal input
rlabel metal2 s 83830 0 83886 800 6 la_data_in[58]
port 199 nsew signal input
rlabel metal2 s 84750 0 84806 800 6 la_data_in[59]
port 200 nsew signal input
rlabel metal2 s 36266 0 36322 800 6 la_data_in[5]
port 201 nsew signal input
rlabel metal2 s 85578 0 85634 800 6 la_data_in[60]
port 202 nsew signal input
rlabel metal2 s 86498 0 86554 800 6 la_data_in[61]
port 203 nsew signal input
rlabel metal2 s 87418 0 87474 800 6 la_data_in[62]
port 204 nsew signal input
rlabel metal2 s 88338 0 88394 800 6 la_data_in[63]
port 205 nsew signal input
rlabel metal2 s 89166 0 89222 800 6 la_data_in[64]
port 206 nsew signal input
rlabel metal2 s 90086 0 90142 800 6 la_data_in[65]
port 207 nsew signal input
rlabel metal2 s 91006 0 91062 800 6 la_data_in[66]
port 208 nsew signal input
rlabel metal2 s 91926 0 91982 800 6 la_data_in[67]
port 209 nsew signal input
rlabel metal2 s 92754 0 92810 800 6 la_data_in[68]
port 210 nsew signal input
rlabel metal2 s 93674 0 93730 800 6 la_data_in[69]
port 211 nsew signal input
rlabel metal2 s 37186 0 37242 800 6 la_data_in[6]
port 212 nsew signal input
rlabel metal2 s 94594 0 94650 800 6 la_data_in[70]
port 213 nsew signal input
rlabel metal2 s 95514 0 95570 800 6 la_data_in[71]
port 214 nsew signal input
rlabel metal2 s 96342 0 96398 800 6 la_data_in[72]
port 215 nsew signal input
rlabel metal2 s 97262 0 97318 800 6 la_data_in[73]
port 216 nsew signal input
rlabel metal2 s 98182 0 98238 800 6 la_data_in[74]
port 217 nsew signal input
rlabel metal2 s 99102 0 99158 800 6 la_data_in[75]
port 218 nsew signal input
rlabel metal2 s 100022 0 100078 800 6 la_data_in[76]
port 219 nsew signal input
rlabel metal2 s 100850 0 100906 800 6 la_data_in[77]
port 220 nsew signal input
rlabel metal2 s 101770 0 101826 800 6 la_data_in[78]
port 221 nsew signal input
rlabel metal2 s 102690 0 102746 800 6 la_data_in[79]
port 222 nsew signal input
rlabel metal2 s 38014 0 38070 800 6 la_data_in[7]
port 223 nsew signal input
rlabel metal2 s 103610 0 103666 800 6 la_data_in[80]
port 224 nsew signal input
rlabel metal2 s 104438 0 104494 800 6 la_data_in[81]
port 225 nsew signal input
rlabel metal2 s 105358 0 105414 800 6 la_data_in[82]
port 226 nsew signal input
rlabel metal2 s 106278 0 106334 800 6 la_data_in[83]
port 227 nsew signal input
rlabel metal2 s 107198 0 107254 800 6 la_data_in[84]
port 228 nsew signal input
rlabel metal2 s 108026 0 108082 800 6 la_data_in[85]
port 229 nsew signal input
rlabel metal2 s 108946 0 109002 800 6 la_data_in[86]
port 230 nsew signal input
rlabel metal2 s 109866 0 109922 800 6 la_data_in[87]
port 231 nsew signal input
rlabel metal2 s 110786 0 110842 800 6 la_data_in[88]
port 232 nsew signal input
rlabel metal2 s 111614 0 111670 800 6 la_data_in[89]
port 233 nsew signal input
rlabel metal2 s 38934 0 38990 800 6 la_data_in[8]
port 234 nsew signal input
rlabel metal2 s 112534 0 112590 800 6 la_data_in[90]
port 235 nsew signal input
rlabel metal2 s 113454 0 113510 800 6 la_data_in[91]
port 236 nsew signal input
rlabel metal2 s 114374 0 114430 800 6 la_data_in[92]
port 237 nsew signal input
rlabel metal2 s 115202 0 115258 800 6 la_data_in[93]
port 238 nsew signal input
rlabel metal2 s 116122 0 116178 800 6 la_data_in[94]
port 239 nsew signal input
rlabel metal2 s 117042 0 117098 800 6 la_data_in[95]
port 240 nsew signal input
rlabel metal2 s 117962 0 118018 800 6 la_data_in[96]
port 241 nsew signal input
rlabel metal2 s 118790 0 118846 800 6 la_data_in[97]
port 242 nsew signal input
rlabel metal2 s 119710 0 119766 800 6 la_data_in[98]
port 243 nsew signal input
rlabel metal2 s 120630 0 120686 800 6 la_data_in[99]
port 244 nsew signal input
rlabel metal2 s 39854 0 39910 800 6 la_data_in[9]
port 245 nsew signal input
rlabel metal2 s 32034 0 32090 800 6 la_data_out[0]
port 246 nsew signal output
rlabel metal2 s 121826 0 121882 800 6 la_data_out[100]
port 247 nsew signal output
rlabel metal2 s 122746 0 122802 800 6 la_data_out[101]
port 248 nsew signal output
rlabel metal2 s 123574 0 123630 800 6 la_data_out[102]
port 249 nsew signal output
rlabel metal2 s 124494 0 124550 800 6 la_data_out[103]
port 250 nsew signal output
rlabel metal2 s 125414 0 125470 800 6 la_data_out[104]
port 251 nsew signal output
rlabel metal2 s 126334 0 126390 800 6 la_data_out[105]
port 252 nsew signal output
rlabel metal2 s 127162 0 127218 800 6 la_data_out[106]
port 253 nsew signal output
rlabel metal2 s 128082 0 128138 800 6 la_data_out[107]
port 254 nsew signal output
rlabel metal2 s 129002 0 129058 800 6 la_data_out[108]
port 255 nsew signal output
rlabel metal2 s 129922 0 129978 800 6 la_data_out[109]
port 256 nsew signal output
rlabel metal2 s 41050 0 41106 800 6 la_data_out[10]
port 257 nsew signal output
rlabel metal2 s 130750 0 130806 800 6 la_data_out[110]
port 258 nsew signal output
rlabel metal2 s 131670 0 131726 800 6 la_data_out[111]
port 259 nsew signal output
rlabel metal2 s 132590 0 132646 800 6 la_data_out[112]
port 260 nsew signal output
rlabel metal2 s 133510 0 133566 800 6 la_data_out[113]
port 261 nsew signal output
rlabel metal2 s 134338 0 134394 800 6 la_data_out[114]
port 262 nsew signal output
rlabel metal2 s 135258 0 135314 800 6 la_data_out[115]
port 263 nsew signal output
rlabel metal2 s 136178 0 136234 800 6 la_data_out[116]
port 264 nsew signal output
rlabel metal2 s 137098 0 137154 800 6 la_data_out[117]
port 265 nsew signal output
rlabel metal2 s 137926 0 137982 800 6 la_data_out[118]
port 266 nsew signal output
rlabel metal2 s 138846 0 138902 800 6 la_data_out[119]
port 267 nsew signal output
rlabel metal2 s 41970 0 42026 800 6 la_data_out[11]
port 268 nsew signal output
rlabel metal2 s 139766 0 139822 800 6 la_data_out[120]
port 269 nsew signal output
rlabel metal2 s 140686 0 140742 800 6 la_data_out[121]
port 270 nsew signal output
rlabel metal2 s 141514 0 141570 800 6 la_data_out[122]
port 271 nsew signal output
rlabel metal2 s 142434 0 142490 800 6 la_data_out[123]
port 272 nsew signal output
rlabel metal2 s 143354 0 143410 800 6 la_data_out[124]
port 273 nsew signal output
rlabel metal2 s 144274 0 144330 800 6 la_data_out[125]
port 274 nsew signal output
rlabel metal2 s 145102 0 145158 800 6 la_data_out[126]
port 275 nsew signal output
rlabel metal2 s 146022 0 146078 800 6 la_data_out[127]
port 276 nsew signal output
rlabel metal2 s 42798 0 42854 800 6 la_data_out[12]
port 277 nsew signal output
rlabel metal2 s 43718 0 43774 800 6 la_data_out[13]
port 278 nsew signal output
rlabel metal2 s 44638 0 44694 800 6 la_data_out[14]
port 279 nsew signal output
rlabel metal2 s 45558 0 45614 800 6 la_data_out[15]
port 280 nsew signal output
rlabel metal2 s 46386 0 46442 800 6 la_data_out[16]
port 281 nsew signal output
rlabel metal2 s 47306 0 47362 800 6 la_data_out[17]
port 282 nsew signal output
rlabel metal2 s 48226 0 48282 800 6 la_data_out[18]
port 283 nsew signal output
rlabel metal2 s 49146 0 49202 800 6 la_data_out[19]
port 284 nsew signal output
rlabel metal2 s 32954 0 33010 800 6 la_data_out[1]
port 285 nsew signal output
rlabel metal2 s 50066 0 50122 800 6 la_data_out[20]
port 286 nsew signal output
rlabel metal2 s 50894 0 50950 800 6 la_data_out[21]
port 287 nsew signal output
rlabel metal2 s 51814 0 51870 800 6 la_data_out[22]
port 288 nsew signal output
rlabel metal2 s 52734 0 52790 800 6 la_data_out[23]
port 289 nsew signal output
rlabel metal2 s 53654 0 53710 800 6 la_data_out[24]
port 290 nsew signal output
rlabel metal2 s 54482 0 54538 800 6 la_data_out[25]
port 291 nsew signal output
rlabel metal2 s 55402 0 55458 800 6 la_data_out[26]
port 292 nsew signal output
rlabel metal2 s 56322 0 56378 800 6 la_data_out[27]
port 293 nsew signal output
rlabel metal2 s 57242 0 57298 800 6 la_data_out[28]
port 294 nsew signal output
rlabel metal2 s 58070 0 58126 800 6 la_data_out[29]
port 295 nsew signal output
rlabel metal2 s 33874 0 33930 800 6 la_data_out[2]
port 296 nsew signal output
rlabel metal2 s 58990 0 59046 800 6 la_data_out[30]
port 297 nsew signal output
rlabel metal2 s 59910 0 59966 800 6 la_data_out[31]
port 298 nsew signal output
rlabel metal2 s 60830 0 60886 800 6 la_data_out[32]
port 299 nsew signal output
rlabel metal2 s 61658 0 61714 800 6 la_data_out[33]
port 300 nsew signal output
rlabel metal2 s 62578 0 62634 800 6 la_data_out[34]
port 301 nsew signal output
rlabel metal2 s 63498 0 63554 800 6 la_data_out[35]
port 302 nsew signal output
rlabel metal2 s 64418 0 64474 800 6 la_data_out[36]
port 303 nsew signal output
rlabel metal2 s 65246 0 65302 800 6 la_data_out[37]
port 304 nsew signal output
rlabel metal2 s 66166 0 66222 800 6 la_data_out[38]
port 305 nsew signal output
rlabel metal2 s 67086 0 67142 800 6 la_data_out[39]
port 306 nsew signal output
rlabel metal2 s 34794 0 34850 800 6 la_data_out[3]
port 307 nsew signal output
rlabel metal2 s 68006 0 68062 800 6 la_data_out[40]
port 308 nsew signal output
rlabel metal2 s 68834 0 68890 800 6 la_data_out[41]
port 309 nsew signal output
rlabel metal2 s 69754 0 69810 800 6 la_data_out[42]
port 310 nsew signal output
rlabel metal2 s 70674 0 70730 800 6 la_data_out[43]
port 311 nsew signal output
rlabel metal2 s 71594 0 71650 800 6 la_data_out[44]
port 312 nsew signal output
rlabel metal2 s 72422 0 72478 800 6 la_data_out[45]
port 313 nsew signal output
rlabel metal2 s 73342 0 73398 800 6 la_data_out[46]
port 314 nsew signal output
rlabel metal2 s 74262 0 74318 800 6 la_data_out[47]
port 315 nsew signal output
rlabel metal2 s 75182 0 75238 800 6 la_data_out[48]
port 316 nsew signal output
rlabel metal2 s 76010 0 76066 800 6 la_data_out[49]
port 317 nsew signal output
rlabel metal2 s 35622 0 35678 800 6 la_data_out[4]
port 318 nsew signal output
rlabel metal2 s 76930 0 76986 800 6 la_data_out[50]
port 319 nsew signal output
rlabel metal2 s 77850 0 77906 800 6 la_data_out[51]
port 320 nsew signal output
rlabel metal2 s 78770 0 78826 800 6 la_data_out[52]
port 321 nsew signal output
rlabel metal2 s 79598 0 79654 800 6 la_data_out[53]
port 322 nsew signal output
rlabel metal2 s 80518 0 80574 800 6 la_data_out[54]
port 323 nsew signal output
rlabel metal2 s 81438 0 81494 800 6 la_data_out[55]
port 324 nsew signal output
rlabel metal2 s 82358 0 82414 800 6 la_data_out[56]
port 325 nsew signal output
rlabel metal2 s 83186 0 83242 800 6 la_data_out[57]
port 326 nsew signal output
rlabel metal2 s 84106 0 84162 800 6 la_data_out[58]
port 327 nsew signal output
rlabel metal2 s 85026 0 85082 800 6 la_data_out[59]
port 328 nsew signal output
rlabel metal2 s 36542 0 36598 800 6 la_data_out[5]
port 329 nsew signal output
rlabel metal2 s 85946 0 86002 800 6 la_data_out[60]
port 330 nsew signal output
rlabel metal2 s 86774 0 86830 800 6 la_data_out[61]
port 331 nsew signal output
rlabel metal2 s 87694 0 87750 800 6 la_data_out[62]
port 332 nsew signal output
rlabel metal2 s 88614 0 88670 800 6 la_data_out[63]
port 333 nsew signal output
rlabel metal2 s 89534 0 89590 800 6 la_data_out[64]
port 334 nsew signal output
rlabel metal2 s 90362 0 90418 800 6 la_data_out[65]
port 335 nsew signal output
rlabel metal2 s 91282 0 91338 800 6 la_data_out[66]
port 336 nsew signal output
rlabel metal2 s 92202 0 92258 800 6 la_data_out[67]
port 337 nsew signal output
rlabel metal2 s 93122 0 93178 800 6 la_data_out[68]
port 338 nsew signal output
rlabel metal2 s 93950 0 94006 800 6 la_data_out[69]
port 339 nsew signal output
rlabel metal2 s 37462 0 37518 800 6 la_data_out[6]
port 340 nsew signal output
rlabel metal2 s 94870 0 94926 800 6 la_data_out[70]
port 341 nsew signal output
rlabel metal2 s 95790 0 95846 800 6 la_data_out[71]
port 342 nsew signal output
rlabel metal2 s 96710 0 96766 800 6 la_data_out[72]
port 343 nsew signal output
rlabel metal2 s 97538 0 97594 800 6 la_data_out[73]
port 344 nsew signal output
rlabel metal2 s 98458 0 98514 800 6 la_data_out[74]
port 345 nsew signal output
rlabel metal2 s 99378 0 99434 800 6 la_data_out[75]
port 346 nsew signal output
rlabel metal2 s 100298 0 100354 800 6 la_data_out[76]
port 347 nsew signal output
rlabel metal2 s 101218 0 101274 800 6 la_data_out[77]
port 348 nsew signal output
rlabel metal2 s 102046 0 102102 800 6 la_data_out[78]
port 349 nsew signal output
rlabel metal2 s 102966 0 103022 800 6 la_data_out[79]
port 350 nsew signal output
rlabel metal2 s 38382 0 38438 800 6 la_data_out[7]
port 351 nsew signal output
rlabel metal2 s 103886 0 103942 800 6 la_data_out[80]
port 352 nsew signal output
rlabel metal2 s 104806 0 104862 800 6 la_data_out[81]
port 353 nsew signal output
rlabel metal2 s 105634 0 105690 800 6 la_data_out[82]
port 354 nsew signal output
rlabel metal2 s 106554 0 106610 800 6 la_data_out[83]
port 355 nsew signal output
rlabel metal2 s 107474 0 107530 800 6 la_data_out[84]
port 356 nsew signal output
rlabel metal2 s 108394 0 108450 800 6 la_data_out[85]
port 357 nsew signal output
rlabel metal2 s 109222 0 109278 800 6 la_data_out[86]
port 358 nsew signal output
rlabel metal2 s 110142 0 110198 800 6 la_data_out[87]
port 359 nsew signal output
rlabel metal2 s 111062 0 111118 800 6 la_data_out[88]
port 360 nsew signal output
rlabel metal2 s 111982 0 112038 800 6 la_data_out[89]
port 361 nsew signal output
rlabel metal2 s 39210 0 39266 800 6 la_data_out[8]
port 362 nsew signal output
rlabel metal2 s 112810 0 112866 800 6 la_data_out[90]
port 363 nsew signal output
rlabel metal2 s 113730 0 113786 800 6 la_data_out[91]
port 364 nsew signal output
rlabel metal2 s 114650 0 114706 800 6 la_data_out[92]
port 365 nsew signal output
rlabel metal2 s 115570 0 115626 800 6 la_data_out[93]
port 366 nsew signal output
rlabel metal2 s 116398 0 116454 800 6 la_data_out[94]
port 367 nsew signal output
rlabel metal2 s 117318 0 117374 800 6 la_data_out[95]
port 368 nsew signal output
rlabel metal2 s 118238 0 118294 800 6 la_data_out[96]
port 369 nsew signal output
rlabel metal2 s 119158 0 119214 800 6 la_data_out[97]
port 370 nsew signal output
rlabel metal2 s 119986 0 120042 800 6 la_data_out[98]
port 371 nsew signal output
rlabel metal2 s 120906 0 120962 800 6 la_data_out[99]
port 372 nsew signal output
rlabel metal2 s 40130 0 40186 800 6 la_data_out[9]
port 373 nsew signal output
rlabel metal2 s 32402 0 32458 800 6 la_oenb[0]
port 374 nsew signal input
rlabel metal2 s 122102 0 122158 800 6 la_oenb[100]
port 375 nsew signal input
rlabel metal2 s 123022 0 123078 800 6 la_oenb[101]
port 376 nsew signal input
rlabel metal2 s 123942 0 123998 800 6 la_oenb[102]
port 377 nsew signal input
rlabel metal2 s 124770 0 124826 800 6 la_oenb[103]
port 378 nsew signal input
rlabel metal2 s 125690 0 125746 800 6 la_oenb[104]
port 379 nsew signal input
rlabel metal2 s 126610 0 126666 800 6 la_oenb[105]
port 380 nsew signal input
rlabel metal2 s 127530 0 127586 800 6 la_oenb[106]
port 381 nsew signal input
rlabel metal2 s 128358 0 128414 800 6 la_oenb[107]
port 382 nsew signal input
rlabel metal2 s 129278 0 129334 800 6 la_oenb[108]
port 383 nsew signal input
rlabel metal2 s 130198 0 130254 800 6 la_oenb[109]
port 384 nsew signal input
rlabel metal2 s 41326 0 41382 800 6 la_oenb[10]
port 385 nsew signal input
rlabel metal2 s 131118 0 131174 800 6 la_oenb[110]
port 386 nsew signal input
rlabel metal2 s 131946 0 132002 800 6 la_oenb[111]
port 387 nsew signal input
rlabel metal2 s 132866 0 132922 800 6 la_oenb[112]
port 388 nsew signal input
rlabel metal2 s 133786 0 133842 800 6 la_oenb[113]
port 389 nsew signal input
rlabel metal2 s 134706 0 134762 800 6 la_oenb[114]
port 390 nsew signal input
rlabel metal2 s 135534 0 135590 800 6 la_oenb[115]
port 391 nsew signal input
rlabel metal2 s 136454 0 136510 800 6 la_oenb[116]
port 392 nsew signal input
rlabel metal2 s 137374 0 137430 800 6 la_oenb[117]
port 393 nsew signal input
rlabel metal2 s 138294 0 138350 800 6 la_oenb[118]
port 394 nsew signal input
rlabel metal2 s 139122 0 139178 800 6 la_oenb[119]
port 395 nsew signal input
rlabel metal2 s 42246 0 42302 800 6 la_oenb[11]
port 396 nsew signal input
rlabel metal2 s 140042 0 140098 800 6 la_oenb[120]
port 397 nsew signal input
rlabel metal2 s 140962 0 141018 800 6 la_oenb[121]
port 398 nsew signal input
rlabel metal2 s 141882 0 141938 800 6 la_oenb[122]
port 399 nsew signal input
rlabel metal2 s 142710 0 142766 800 6 la_oenb[123]
port 400 nsew signal input
rlabel metal2 s 143630 0 143686 800 6 la_oenb[124]
port 401 nsew signal input
rlabel metal2 s 144550 0 144606 800 6 la_oenb[125]
port 402 nsew signal input
rlabel metal2 s 145470 0 145526 800 6 la_oenb[126]
port 403 nsew signal input
rlabel metal2 s 146298 0 146354 800 6 la_oenb[127]
port 404 nsew signal input
rlabel metal2 s 43166 0 43222 800 6 la_oenb[12]
port 405 nsew signal input
rlabel metal2 s 43994 0 44050 800 6 la_oenb[13]
port 406 nsew signal input
rlabel metal2 s 44914 0 44970 800 6 la_oenb[14]
port 407 nsew signal input
rlabel metal2 s 45834 0 45890 800 6 la_oenb[15]
port 408 nsew signal input
rlabel metal2 s 46754 0 46810 800 6 la_oenb[16]
port 409 nsew signal input
rlabel metal2 s 47582 0 47638 800 6 la_oenb[17]
port 410 nsew signal input
rlabel metal2 s 48502 0 48558 800 6 la_oenb[18]
port 411 nsew signal input
rlabel metal2 s 49422 0 49478 800 6 la_oenb[19]
port 412 nsew signal input
rlabel metal2 s 33230 0 33286 800 6 la_oenb[1]
port 413 nsew signal input
rlabel metal2 s 50342 0 50398 800 6 la_oenb[20]
port 414 nsew signal input
rlabel metal2 s 51262 0 51318 800 6 la_oenb[21]
port 415 nsew signal input
rlabel metal2 s 52090 0 52146 800 6 la_oenb[22]
port 416 nsew signal input
rlabel metal2 s 53010 0 53066 800 6 la_oenb[23]
port 417 nsew signal input
rlabel metal2 s 53930 0 53986 800 6 la_oenb[24]
port 418 nsew signal input
rlabel metal2 s 54850 0 54906 800 6 la_oenb[25]
port 419 nsew signal input
rlabel metal2 s 55678 0 55734 800 6 la_oenb[26]
port 420 nsew signal input
rlabel metal2 s 56598 0 56654 800 6 la_oenb[27]
port 421 nsew signal input
rlabel metal2 s 57518 0 57574 800 6 la_oenb[28]
port 422 nsew signal input
rlabel metal2 s 58438 0 58494 800 6 la_oenb[29]
port 423 nsew signal input
rlabel metal2 s 34150 0 34206 800 6 la_oenb[2]
port 424 nsew signal input
rlabel metal2 s 59266 0 59322 800 6 la_oenb[30]
port 425 nsew signal input
rlabel metal2 s 60186 0 60242 800 6 la_oenb[31]
port 426 nsew signal input
rlabel metal2 s 61106 0 61162 800 6 la_oenb[32]
port 427 nsew signal input
rlabel metal2 s 62026 0 62082 800 6 la_oenb[33]
port 428 nsew signal input
rlabel metal2 s 62854 0 62910 800 6 la_oenb[34]
port 429 nsew signal input
rlabel metal2 s 63774 0 63830 800 6 la_oenb[35]
port 430 nsew signal input
rlabel metal2 s 64694 0 64750 800 6 la_oenb[36]
port 431 nsew signal input
rlabel metal2 s 65614 0 65670 800 6 la_oenb[37]
port 432 nsew signal input
rlabel metal2 s 66442 0 66498 800 6 la_oenb[38]
port 433 nsew signal input
rlabel metal2 s 67362 0 67418 800 6 la_oenb[39]
port 434 nsew signal input
rlabel metal2 s 35070 0 35126 800 6 la_oenb[3]
port 435 nsew signal input
rlabel metal2 s 68282 0 68338 800 6 la_oenb[40]
port 436 nsew signal input
rlabel metal2 s 69202 0 69258 800 6 la_oenb[41]
port 437 nsew signal input
rlabel metal2 s 70030 0 70086 800 6 la_oenb[42]
port 438 nsew signal input
rlabel metal2 s 70950 0 71006 800 6 la_oenb[43]
port 439 nsew signal input
rlabel metal2 s 71870 0 71926 800 6 la_oenb[44]
port 440 nsew signal input
rlabel metal2 s 72790 0 72846 800 6 la_oenb[45]
port 441 nsew signal input
rlabel metal2 s 73618 0 73674 800 6 la_oenb[46]
port 442 nsew signal input
rlabel metal2 s 74538 0 74594 800 6 la_oenb[47]
port 443 nsew signal input
rlabel metal2 s 75458 0 75514 800 6 la_oenb[48]
port 444 nsew signal input
rlabel metal2 s 76378 0 76434 800 6 la_oenb[49]
port 445 nsew signal input
rlabel metal2 s 35990 0 36046 800 6 la_oenb[4]
port 446 nsew signal input
rlabel metal2 s 77206 0 77262 800 6 la_oenb[50]
port 447 nsew signal input
rlabel metal2 s 78126 0 78182 800 6 la_oenb[51]
port 448 nsew signal input
rlabel metal2 s 79046 0 79102 800 6 la_oenb[52]
port 449 nsew signal input
rlabel metal2 s 79966 0 80022 800 6 la_oenb[53]
port 450 nsew signal input
rlabel metal2 s 80794 0 80850 800 6 la_oenb[54]
port 451 nsew signal input
rlabel metal2 s 81714 0 81770 800 6 la_oenb[55]
port 452 nsew signal input
rlabel metal2 s 82634 0 82690 800 6 la_oenb[56]
port 453 nsew signal input
rlabel metal2 s 83554 0 83610 800 6 la_oenb[57]
port 454 nsew signal input
rlabel metal2 s 84382 0 84438 800 6 la_oenb[58]
port 455 nsew signal input
rlabel metal2 s 85302 0 85358 800 6 la_oenb[59]
port 456 nsew signal input
rlabel metal2 s 36818 0 36874 800 6 la_oenb[5]
port 457 nsew signal input
rlabel metal2 s 86222 0 86278 800 6 la_oenb[60]
port 458 nsew signal input
rlabel metal2 s 87142 0 87198 800 6 la_oenb[61]
port 459 nsew signal input
rlabel metal2 s 87970 0 88026 800 6 la_oenb[62]
port 460 nsew signal input
rlabel metal2 s 88890 0 88946 800 6 la_oenb[63]
port 461 nsew signal input
rlabel metal2 s 89810 0 89866 800 6 la_oenb[64]
port 462 nsew signal input
rlabel metal2 s 90730 0 90786 800 6 la_oenb[65]
port 463 nsew signal input
rlabel metal2 s 91558 0 91614 800 6 la_oenb[66]
port 464 nsew signal input
rlabel metal2 s 92478 0 92534 800 6 la_oenb[67]
port 465 nsew signal input
rlabel metal2 s 93398 0 93454 800 6 la_oenb[68]
port 466 nsew signal input
rlabel metal2 s 94318 0 94374 800 6 la_oenb[69]
port 467 nsew signal input
rlabel metal2 s 37738 0 37794 800 6 la_oenb[6]
port 468 nsew signal input
rlabel metal2 s 95146 0 95202 800 6 la_oenb[70]
port 469 nsew signal input
rlabel metal2 s 96066 0 96122 800 6 la_oenb[71]
port 470 nsew signal input
rlabel metal2 s 96986 0 97042 800 6 la_oenb[72]
port 471 nsew signal input
rlabel metal2 s 97906 0 97962 800 6 la_oenb[73]
port 472 nsew signal input
rlabel metal2 s 98826 0 98882 800 6 la_oenb[74]
port 473 nsew signal input
rlabel metal2 s 99654 0 99710 800 6 la_oenb[75]
port 474 nsew signal input
rlabel metal2 s 100574 0 100630 800 6 la_oenb[76]
port 475 nsew signal input
rlabel metal2 s 101494 0 101550 800 6 la_oenb[77]
port 476 nsew signal input
rlabel metal2 s 102414 0 102470 800 6 la_oenb[78]
port 477 nsew signal input
rlabel metal2 s 103242 0 103298 800 6 la_oenb[79]
port 478 nsew signal input
rlabel metal2 s 38658 0 38714 800 6 la_oenb[7]
port 479 nsew signal input
rlabel metal2 s 104162 0 104218 800 6 la_oenb[80]
port 480 nsew signal input
rlabel metal2 s 105082 0 105138 800 6 la_oenb[81]
port 481 nsew signal input
rlabel metal2 s 106002 0 106058 800 6 la_oenb[82]
port 482 nsew signal input
rlabel metal2 s 106830 0 106886 800 6 la_oenb[83]
port 483 nsew signal input
rlabel metal2 s 107750 0 107806 800 6 la_oenb[84]
port 484 nsew signal input
rlabel metal2 s 108670 0 108726 800 6 la_oenb[85]
port 485 nsew signal input
rlabel metal2 s 109590 0 109646 800 6 la_oenb[86]
port 486 nsew signal input
rlabel metal2 s 110418 0 110474 800 6 la_oenb[87]
port 487 nsew signal input
rlabel metal2 s 111338 0 111394 800 6 la_oenb[88]
port 488 nsew signal input
rlabel metal2 s 112258 0 112314 800 6 la_oenb[89]
port 489 nsew signal input
rlabel metal2 s 39578 0 39634 800 6 la_oenb[8]
port 490 nsew signal input
rlabel metal2 s 113178 0 113234 800 6 la_oenb[90]
port 491 nsew signal input
rlabel metal2 s 114006 0 114062 800 6 la_oenb[91]
port 492 nsew signal input
rlabel metal2 s 114926 0 114982 800 6 la_oenb[92]
port 493 nsew signal input
rlabel metal2 s 115846 0 115902 800 6 la_oenb[93]
port 494 nsew signal input
rlabel metal2 s 116766 0 116822 800 6 la_oenb[94]
port 495 nsew signal input
rlabel metal2 s 117594 0 117650 800 6 la_oenb[95]
port 496 nsew signal input
rlabel metal2 s 118514 0 118570 800 6 la_oenb[96]
port 497 nsew signal input
rlabel metal2 s 119434 0 119490 800 6 la_oenb[97]
port 498 nsew signal input
rlabel metal2 s 120354 0 120410 800 6 la_oenb[98]
port 499 nsew signal input
rlabel metal2 s 121182 0 121238 800 6 la_oenb[99]
port 500 nsew signal input
rlabel metal2 s 40406 0 40462 800 6 la_oenb[9]
port 501 nsew signal input
rlabel metal4 s 4208 2128 4528 147472 6 vccd1
port 502 nsew power input
rlabel metal4 s 34928 2128 35248 147472 6 vccd1
port 502 nsew power input
rlabel metal4 s 65648 2128 65968 147472 6 vccd1
port 502 nsew power input
rlabel metal4 s 96368 2128 96688 147472 6 vccd1
port 502 nsew power input
rlabel metal4 s 127088 2128 127408 147472 6 vccd1
port 502 nsew power input
rlabel metal4 s 19568 2128 19888 147472 6 vssd1
port 503 nsew ground input
rlabel metal4 s 50288 2128 50608 147472 6 vssd1
port 503 nsew ground input
rlabel metal4 s 81008 2128 81328 147472 6 vssd1
port 503 nsew ground input
rlabel metal4 s 111728 2128 112048 147472 6 vssd1
port 503 nsew ground input
rlabel metal4 s 142448 2128 142768 147472 6 vssd1
port 503 nsew ground input
rlabel metal2 s 110 0 166 800 6 wb_clk_i
port 504 nsew signal input
rlabel metal2 s 386 0 442 800 6 wb_rst_i
port 505 nsew signal input
rlabel metal2 s 662 0 718 800 6 wbs_ack_o
port 506 nsew signal output
rlabel metal2 s 1858 0 1914 800 6 wbs_adr_i[0]
port 507 nsew signal input
rlabel metal2 s 12070 0 12126 800 6 wbs_adr_i[10]
port 508 nsew signal input
rlabel metal2 s 12898 0 12954 800 6 wbs_adr_i[11]
port 509 nsew signal input
rlabel metal2 s 13818 0 13874 800 6 wbs_adr_i[12]
port 510 nsew signal input
rlabel metal2 s 14738 0 14794 800 6 wbs_adr_i[13]
port 511 nsew signal input
rlabel metal2 s 15658 0 15714 800 6 wbs_adr_i[14]
port 512 nsew signal input
rlabel metal2 s 16486 0 16542 800 6 wbs_adr_i[15]
port 513 nsew signal input
rlabel metal2 s 17406 0 17462 800 6 wbs_adr_i[16]
port 514 nsew signal input
rlabel metal2 s 18326 0 18382 800 6 wbs_adr_i[17]
port 515 nsew signal input
rlabel metal2 s 19246 0 19302 800 6 wbs_adr_i[18]
port 516 nsew signal input
rlabel metal2 s 20074 0 20130 800 6 wbs_adr_i[19]
port 517 nsew signal input
rlabel metal2 s 3054 0 3110 800 6 wbs_adr_i[1]
port 518 nsew signal input
rlabel metal2 s 20994 0 21050 800 6 wbs_adr_i[20]
port 519 nsew signal input
rlabel metal2 s 21914 0 21970 800 6 wbs_adr_i[21]
port 520 nsew signal input
rlabel metal2 s 22834 0 22890 800 6 wbs_adr_i[22]
port 521 nsew signal input
rlabel metal2 s 23662 0 23718 800 6 wbs_adr_i[23]
port 522 nsew signal input
rlabel metal2 s 24582 0 24638 800 6 wbs_adr_i[24]
port 523 nsew signal input
rlabel metal2 s 25502 0 25558 800 6 wbs_adr_i[25]
port 524 nsew signal input
rlabel metal2 s 26422 0 26478 800 6 wbs_adr_i[26]
port 525 nsew signal input
rlabel metal2 s 27250 0 27306 800 6 wbs_adr_i[27]
port 526 nsew signal input
rlabel metal2 s 28170 0 28226 800 6 wbs_adr_i[28]
port 527 nsew signal input
rlabel metal2 s 29090 0 29146 800 6 wbs_adr_i[29]
port 528 nsew signal input
rlabel metal2 s 4250 0 4306 800 6 wbs_adr_i[2]
port 529 nsew signal input
rlabel metal2 s 30010 0 30066 800 6 wbs_adr_i[30]
port 530 nsew signal input
rlabel metal2 s 30838 0 30894 800 6 wbs_adr_i[31]
port 531 nsew signal input
rlabel metal2 s 5446 0 5502 800 6 wbs_adr_i[3]
port 532 nsew signal input
rlabel metal2 s 6642 0 6698 800 6 wbs_adr_i[4]
port 533 nsew signal input
rlabel metal2 s 7562 0 7618 800 6 wbs_adr_i[5]
port 534 nsew signal input
rlabel metal2 s 8482 0 8538 800 6 wbs_adr_i[6]
port 535 nsew signal input
rlabel metal2 s 9310 0 9366 800 6 wbs_adr_i[7]
port 536 nsew signal input
rlabel metal2 s 10230 0 10286 800 6 wbs_adr_i[8]
port 537 nsew signal input
rlabel metal2 s 11150 0 11206 800 6 wbs_adr_i[9]
port 538 nsew signal input
rlabel metal2 s 938 0 994 800 6 wbs_cyc_i
port 539 nsew signal input
rlabel metal2 s 2134 0 2190 800 6 wbs_dat_i[0]
port 540 nsew signal input
rlabel metal2 s 12346 0 12402 800 6 wbs_dat_i[10]
port 541 nsew signal input
rlabel metal2 s 13266 0 13322 800 6 wbs_dat_i[11]
port 542 nsew signal input
rlabel metal2 s 14094 0 14150 800 6 wbs_dat_i[12]
port 543 nsew signal input
rlabel metal2 s 15014 0 15070 800 6 wbs_dat_i[13]
port 544 nsew signal input
rlabel metal2 s 15934 0 15990 800 6 wbs_dat_i[14]
port 545 nsew signal input
rlabel metal2 s 16854 0 16910 800 6 wbs_dat_i[15]
port 546 nsew signal input
rlabel metal2 s 17682 0 17738 800 6 wbs_dat_i[16]
port 547 nsew signal input
rlabel metal2 s 18602 0 18658 800 6 wbs_dat_i[17]
port 548 nsew signal input
rlabel metal2 s 19522 0 19578 800 6 wbs_dat_i[18]
port 549 nsew signal input
rlabel metal2 s 20442 0 20498 800 6 wbs_dat_i[19]
port 550 nsew signal input
rlabel metal2 s 3330 0 3386 800 6 wbs_dat_i[1]
port 551 nsew signal input
rlabel metal2 s 21270 0 21326 800 6 wbs_dat_i[20]
port 552 nsew signal input
rlabel metal2 s 22190 0 22246 800 6 wbs_dat_i[21]
port 553 nsew signal input
rlabel metal2 s 23110 0 23166 800 6 wbs_dat_i[22]
port 554 nsew signal input
rlabel metal2 s 24030 0 24086 800 6 wbs_dat_i[23]
port 555 nsew signal input
rlabel metal2 s 24858 0 24914 800 6 wbs_dat_i[24]
port 556 nsew signal input
rlabel metal2 s 25778 0 25834 800 6 wbs_dat_i[25]
port 557 nsew signal input
rlabel metal2 s 26698 0 26754 800 6 wbs_dat_i[26]
port 558 nsew signal input
rlabel metal2 s 27618 0 27674 800 6 wbs_dat_i[27]
port 559 nsew signal input
rlabel metal2 s 28446 0 28502 800 6 wbs_dat_i[28]
port 560 nsew signal input
rlabel metal2 s 29366 0 29422 800 6 wbs_dat_i[29]
port 561 nsew signal input
rlabel metal2 s 4526 0 4582 800 6 wbs_dat_i[2]
port 562 nsew signal input
rlabel metal2 s 30286 0 30342 800 6 wbs_dat_i[30]
port 563 nsew signal input
rlabel metal2 s 31206 0 31262 800 6 wbs_dat_i[31]
port 564 nsew signal input
rlabel metal2 s 5722 0 5778 800 6 wbs_dat_i[3]
port 565 nsew signal input
rlabel metal2 s 6918 0 6974 800 6 wbs_dat_i[4]
port 566 nsew signal input
rlabel metal2 s 7838 0 7894 800 6 wbs_dat_i[5]
port 567 nsew signal input
rlabel metal2 s 8758 0 8814 800 6 wbs_dat_i[6]
port 568 nsew signal input
rlabel metal2 s 9678 0 9734 800 6 wbs_dat_i[7]
port 569 nsew signal input
rlabel metal2 s 10506 0 10562 800 6 wbs_dat_i[8]
port 570 nsew signal input
rlabel metal2 s 11426 0 11482 800 6 wbs_dat_i[9]
port 571 nsew signal input
rlabel metal2 s 2502 0 2558 800 6 wbs_dat_o[0]
port 572 nsew signal output
rlabel metal2 s 12622 0 12678 800 6 wbs_dat_o[10]
port 573 nsew signal output
rlabel metal2 s 13542 0 13598 800 6 wbs_dat_o[11]
port 574 nsew signal output
rlabel metal2 s 14462 0 14518 800 6 wbs_dat_o[12]
port 575 nsew signal output
rlabel metal2 s 15290 0 15346 800 6 wbs_dat_o[13]
port 576 nsew signal output
rlabel metal2 s 16210 0 16266 800 6 wbs_dat_o[14]
port 577 nsew signal output
rlabel metal2 s 17130 0 17186 800 6 wbs_dat_o[15]
port 578 nsew signal output
rlabel metal2 s 18050 0 18106 800 6 wbs_dat_o[16]
port 579 nsew signal output
rlabel metal2 s 18878 0 18934 800 6 wbs_dat_o[17]
port 580 nsew signal output
rlabel metal2 s 19798 0 19854 800 6 wbs_dat_o[18]
port 581 nsew signal output
rlabel metal2 s 20718 0 20774 800 6 wbs_dat_o[19]
port 582 nsew signal output
rlabel metal2 s 3698 0 3754 800 6 wbs_dat_o[1]
port 583 nsew signal output
rlabel metal2 s 21638 0 21694 800 6 wbs_dat_o[20]
port 584 nsew signal output
rlabel metal2 s 22466 0 22522 800 6 wbs_dat_o[21]
port 585 nsew signal output
rlabel metal2 s 23386 0 23442 800 6 wbs_dat_o[22]
port 586 nsew signal output
rlabel metal2 s 24306 0 24362 800 6 wbs_dat_o[23]
port 587 nsew signal output
rlabel metal2 s 25226 0 25282 800 6 wbs_dat_o[24]
port 588 nsew signal output
rlabel metal2 s 26054 0 26110 800 6 wbs_dat_o[25]
port 589 nsew signal output
rlabel metal2 s 26974 0 27030 800 6 wbs_dat_o[26]
port 590 nsew signal output
rlabel metal2 s 27894 0 27950 800 6 wbs_dat_o[27]
port 591 nsew signal output
rlabel metal2 s 28814 0 28870 800 6 wbs_dat_o[28]
port 592 nsew signal output
rlabel metal2 s 29642 0 29698 800 6 wbs_dat_o[29]
port 593 nsew signal output
rlabel metal2 s 4894 0 4950 800 6 wbs_dat_o[2]
port 594 nsew signal output
rlabel metal2 s 30562 0 30618 800 6 wbs_dat_o[30]
port 595 nsew signal output
rlabel metal2 s 31482 0 31538 800 6 wbs_dat_o[31]
port 596 nsew signal output
rlabel metal2 s 6090 0 6146 800 6 wbs_dat_o[3]
port 597 nsew signal output
rlabel metal2 s 7286 0 7342 800 6 wbs_dat_o[4]
port 598 nsew signal output
rlabel metal2 s 8114 0 8170 800 6 wbs_dat_o[5]
port 599 nsew signal output
rlabel metal2 s 9034 0 9090 800 6 wbs_dat_o[6]
port 600 nsew signal output
rlabel metal2 s 9954 0 10010 800 6 wbs_dat_o[7]
port 601 nsew signal output
rlabel metal2 s 10874 0 10930 800 6 wbs_dat_o[8]
port 602 nsew signal output
rlabel metal2 s 11702 0 11758 800 6 wbs_dat_o[9]
port 603 nsew signal output
rlabel metal2 s 2778 0 2834 800 6 wbs_sel_i[0]
port 604 nsew signal input
rlabel metal2 s 3974 0 4030 800 6 wbs_sel_i[1]
port 605 nsew signal input
rlabel metal2 s 5170 0 5226 800 6 wbs_sel_i[2]
port 606 nsew signal input
rlabel metal2 s 6366 0 6422 800 6 wbs_sel_i[3]
port 607 nsew signal input
rlabel metal2 s 1306 0 1362 800 6 wbs_stb_i
port 608 nsew signal input
rlabel metal2 s 1582 0 1638 800 6 wbs_we_i
port 609 nsew signal input
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 147459 149603
string LEFview TRUE
string GDS_FILE /project/openlane/user_proj_example/runs/user_proj_example/results/magic/user_proj_example.gds
string GDS_END 57256346
string GDS_START 621000
<< end >>

