`timescale 1ns / 100ps

module sbox2(
    input [5:0] i_data,
    output reg [3:0] o_data
);



    always@(i_data) begin
        case(i_data)
            6'b000000: o_data = 4'b1111; // (0, 0) = 15
            6'b000001: o_data = 4'b0011; // (0, 1) = 3
            6'b000010: o_data = 4'b0001; // (1, 0) = 1
            6'b000011: o_data = 4'b1101; // (1, 1) = 13
            6'b000100: o_data = 4'b1000; // (2, 0) = 8
            6'b000101: o_data = 4'b0100; // (2, 1) = 4
            6'b000110: o_data = 4'b1110; // (3, 0) = 14
            6'b000111: o_data = 4'b0111; // (3, 1) = 7
            6'b001000: o_data = 4'b0110; // (4, 0) = 6
            6'b001001: o_data = 4'b1111; // (4, 1) = 15
            6'b001010: o_data = 4'b1011; // (5, 0) = 11
            6'b001011: o_data = 4'b0010; // (5, 1) = 2
            6'b001100: o_data = 4'b0011; // (6, 0) = 3
            6'b001101: o_data = 4'b1000; // (6, 1) = 8
            6'b001110: o_data = 4'b0100; // (7, 0) = 4
            6'b001111: o_data = 4'b1110; // (7, 1) = 14
            6'b010000: o_data = 4'b1001; // (8, 0) = 9
            6'b010001: o_data = 4'b1100; // (8, 1) = 12
            6'b010010: o_data = 4'b0111; // (9, 0) = 7
            6'b010011: o_data = 4'b0000; // (9, 1) = 0
            6'b010100: o_data = 4'b0010; // (10, 0) = 2
            6'b010101: o_data = 4'b0001; // (10, 1) = 1
            6'b010110: o_data = 4'b1101; // (11, 0) = 13
            6'b010111: o_data = 4'b1010; // (11, 1) = 10
            6'b011000: o_data = 4'b1100; // (12, 0) = 12
            6'b011001: o_data = 4'b0110; // (12, 1) = 6
            6'b011010: o_data = 4'b0000; // (13, 0) = 0
            6'b011011: o_data = 4'b1001; // (13, 1) = 9
            6'b011100: o_data = 4'b0101; // (14, 0) = 5
            6'b011101: o_data = 4'b1011; // (14, 1) = 11
            6'b011110: o_data = 4'b1010; // (15, 0) = 10
            6'b011111: o_data = 4'b0101; // (15, 1) = 5
            6'b100000: o_data = 4'b0000; // (0, 2) = 0
            6'b100001: o_data = 4'b1101; // (0, 3) = 13
            6'b100010: o_data = 4'b1110; // (1, 2) = 14
            6'b100011: o_data = 4'b1000; // (1, 3) = 8
            6'b100100: o_data = 4'b0111; // (2, 2) = 7
            6'b100101: o_data = 4'b1010; // (2, 3) = 10
            6'b100110: o_data = 4'b1011; // (3, 2) = 11
            6'b100111: o_data = 4'b0001; // (3, 3) = 1
            6'b101000: o_data = 4'b1010; // (4, 2) = 10
            6'b101001: o_data = 4'b0011; // (4, 3) = 3
            6'b101010: o_data = 4'b0100; // (5, 2) = 4
            6'b101011: o_data = 4'b1111; // (5, 3) = 15
            6'b101100: o_data = 4'b1101; // (6, 2) = 13
            6'b101101: o_data = 4'b0100; // (6, 3) = 4
            6'b101110: o_data = 4'b0001; // (7, 2) = 1
            6'b101111: o_data = 4'b0010; // (7, 3) = 2
            6'b110000: o_data = 4'b0101; // (8, 2) = 5
            6'b110001: o_data = 4'b1011; // (8, 3) = 11
            6'b110010: o_data = 4'b1000; // (9, 2) = 8
            6'b110011: o_data = 4'b0110; // (9, 3) = 6
            6'b110100: o_data = 4'b1100; // (10, 2) = 12
            6'b110101: o_data = 4'b0111; // (10, 3) = 7
            6'b110110: o_data = 4'b0110; // (11, 2) = 6
            6'b110111: o_data = 4'b1100; // (11, 3) = 12
            6'b111000: o_data = 4'b1001; // (12, 2) = 9
            6'b111001: o_data = 4'b0000; // (12, 3) = 0
            6'b111010: o_data = 4'b0011; // (13, 2) = 3
            6'b111011: o_data = 4'b0101; // (13, 3) = 5
            6'b111100: o_data = 4'b0010; // (14, 2) = 2
            6'b111101: o_data = 4'b1110; // (14, 3) = 14
            6'b111110: o_data = 4'b1111; // (15, 2) = 15
            6'b111111: o_data = 4'b1001; // (15, 3) = 9
        endcase
    end
endmodule
